module memory #(
    parameter SAMPLE_WIDTH = 18,
    parameter ADDR_WIDTH   = 10
)(
    input  wire clk,
    input  wire [ADDR_WIDTH-1:0] addr_a,
        output reg  [SAMPLE_WIDTH-1:0] data_out_a,
        input  wire [ADDR_WIDTH-1:0] addr_b,
        output reg  [SAMPLE_WIDTH-1:0] data_out_b
    );

    (* ram_style = "block" *) reg [SAMPLE_WIDTH-1:0] mem [0:1023];// 1024 samples total

    
    initial begin

    mem[0] = { 8'd57, 8'd59, 2'd0 }; // Age: 57, HR: 159, Class: 0
mem[1] = { 8'd53, 8'd30, 2'd0 }; // Age: 53, HR: 130, Class: 0
mem[2] = { 8'd62, 8'd38, 2'd1 }; // Age: 62, HR: 138, Class: 1
mem[3] = { 8'd61, 8'd38, 2'd1 }; // Age: 61, HR: 138, Class: 1
mem[4] = { 8'd59, 8'd62, 2'd2 }; // Age: 59, HR: 162, Class: 2
mem[5] = { 8'd67, 8'd63, 2'd3 }; // Age: 67, HR: 163, Class: 3
mem[6] = { 8'd64, 8'd40, 2'd3 }; // Age: 64, HR: 140, Class: 3
mem[7] = { 8'd64, 8'd44, 2'd0 }; // Age: 64, HR: 144, Class: 0
mem[8] = { 8'd46, 8'd33, 2'd1 }; // Age: 46, HR: 133, Class: 1
mem[9] = { 8'd63, 8'd54, 2'd3 }; // Age: 63, HR: 154, Class: 3
mem[10] = { 8'd55, 8'd40, 2'd0 }; // Age: 55, HR: 140, Class: 0
mem[11] = { 8'd52, 8'd60, 2'd1 }; // Age: 52, HR: 160, Class: 1
mem[12] = { 8'd38, 8'd29, 2'd0 }; // Age: 38, HR: 129, Class: 0
mem[13] = { 8'd55, 8'd60, 2'd0 }; // Age: 55, HR: 160, Class: 0
mem[14] = { 8'd53, 8'd15, 2'd0 }; // Age: 53, HR: 115, Class: 0
mem[15] = { 8'd44, 8'd35, 2'd0 }; // Age: 44, HR: 135, Class: 0
mem[16] = { 8'd48, 8'd86, 2'd0 }; // Age: 48, HR: 186, Class: 0
mem[17] = { 8'd57, 8'd254, 2'd2 }; // Age: 57, HR: 98, Class: 2
mem[18] = { 8'd54, 8'd47, 2'd0 }; // Age: 54, HR: 147, Class: 0
mem[19] = { 8'd57, 8'd20, 2'd2 }; // Age: 57, HR: 120, Class: 2
mem[20] = { 8'd32, 8'd65, 2'd0 }; // Age: 32, HR: 165, Class: 0
mem[21] = { 8'd56, 8'd23, 2'd3 }; // Age: 56, HR: 123, Class: 3
mem[22] = { 8'd40, 8'd50, 2'd0 }; // Age: 40, HR: 150, Class: 0
mem[23] = { 8'd33, 8'd50, 2'd1 }; // Age: 33, HR: 150, Class: 1
mem[24] = { 8'd50, 8'd60, 2'd0 }; // Age: 50, HR: 160, Class: 0
mem[25] = { 8'd59, 8'd17, 2'd1 }; // Age: 59, HR: 117, Class: 1
mem[26] = { 8'd46, 8'd40, 2'd0 }; // Age: 46, HR: 140, Class: 0
mem[27] = { 8'd51, 8'd22, 2'd3 }; // Age: 51, HR: 122, Class: 3
mem[28] = { 8'd66, 8'd52, 2'd0 }; // Age: 66, HR: 152, Class: 0
mem[29] = { 8'd46, 8'd56, 2'd0 }; // Age: 46, HR: 156, Class: 0
mem[30] = { 8'd55, 8'd55, 2'd0 }; // Age: 55, HR: 155, Class: 0
mem[31] = { 8'd34, 8'd68, 2'd0 }; // Age: 34, HR: 168, Class: 0
mem[32] = { 8'd58, 8'd62, 2'd0 }; // Age: 58, HR: 162, Class: 0
mem[33] = { 8'd64, 8'd5, 2'd0 }; // Age: 64, HR: 105, Class: 0
mem[34] = { 8'd52, 8'd10, 2'd2 }; // Age: 52, HR: 110, Class: 2
mem[35] = { 8'd68, 8'd51, 2'd0 }; // Age: 68, HR: 151, Class: 0
mem[36] = { 8'd49, 8'd20, 2'd1 }; // Age: 49, HR: 120, Class: 1
mem[37] = { 8'd57, 8'd26, 2'd0 }; // Age: 57, HR: 126, Class: 0
mem[38] = { 8'd54, 8'd52, 2'd0 }; // Age: 54, HR: 152, Class: 0
mem[39] = { 8'd48, 8'd3, 2'd1 }; // Age: 48, HR: 103, Class: 1
mem[40] = { 8'd61, 8'd13, 2'd1 }; // Age: 61, HR: 113, Class: 1
mem[41] = { 8'd57, 8'd40, 2'd0 }; // Age: 57, HR: 140, Class: 0
mem[42] = { 8'd63, 8'd254, 2'd1 }; // Age: 63, HR: 98, Class: 1
mem[43] = { 8'd58, 8'd225, 2'd0 }; // Age: 58, HR: 69, Class: 0
mem[44] = { 8'd69, 8'd46, 2'd2 }; // Age: 69, HR: 146, Class: 2
mem[45] = { 8'd61, 8'd17, 2'd2 }; // Age: 61, HR: 117, Class: 2
mem[46] = { 8'd51, 8'd50, 2'd1 }; // Age: 51, HR: 150, Class: 1
mem[47] = { 8'd52, 8'd238, 2'd1 }; // Age: 52, HR: 82, Class: 1
mem[48] = { 8'd61, 8'd45, 2'd2 }; // Age: 61, HR: 145, Class: 2
mem[49] = { 8'd55, 8'd10, 2'd1 }; // Age: 55, HR: 110, Class: 1
mem[50] = { 8'd46, 8'd24, 2'd1 }; // Age: 46, HR: 124, Class: 1
mem[51] = { 8'd54, 8'd47, 2'd0 }; // Age: 54, HR: 147, Class: 0
mem[52] = { 8'd59, 8'd40, 2'd0 }; // Age: 59, HR: 140, Class: 0
mem[53] = { 8'd61, 8'd0, 2'd3 }; // Age: 61, HR: 100, Class: 3
mem[54] = { 8'd54, 8'd50, 2'd1 }; // Age: 54, HR: 150, Class: 1
mem[55] = { 8'd64, 8'd44, 2'd0 }; // Age: 64, HR: 144, Class: 0
mem[56] = { 8'd53, 8'd22, 2'd1 }; // Age: 53, HR: 122, Class: 1
mem[57] = { 8'd52, 8'd69, 2'd0 }; // Age: 52, HR: 169, Class: 0
mem[58] = { 8'd71, 8'd25, 2'd0 }; // Age: 71, HR: 125, Class: 0
mem[59] = { 8'd46, 8'd20, 2'd0 }; // Age: 46, HR: 120, Class: 0
mem[60] = { 8'd38, 8'd66, 2'd2 }; // Age: 38, HR: 166, Class: 2
mem[61] = { 8'd35, 8'd85, 2'd0 }; // Age: 35, HR: 185, Class: 0
mem[62] = { 8'd44, 8'd73, 2'd0 }; // Age: 44, HR: 173, Class: 0
mem[63] = { 8'd41, 8'd63, 2'd0 }; // Age: 41, HR: 163, Class: 0
mem[64] = { 8'd54, 8'd40, 2'd3 }; // Age: 54, HR: 140, Class: 3
mem[65] = { 8'd40, 8'd38, 2'd0 }; // Age: 40, HR: 138, Class: 0
mem[66] = { 8'd52, 8'd10, 2'd1 }; // Age: 52, HR: 110, Class: 1
mem[67] = { 8'd39, 8'd70, 2'd0 }; // Age: 39, HR: 170, Class: 0
mem[68] = { 8'd62, 8'd45, 2'd3 }; // Age: 62, HR: 145, Class: 3
mem[69] = { 8'd43, 8'd18, 2'd0 }; // Age: 43, HR: 118, Class: 0
mem[70] = { 8'd54, 8'd75, 2'd0 }; // Age: 54, HR: 175, Class: 0
mem[71] = { 8'd52, 8'd39, 2'd0 }; // Age: 52, HR: 139, Class: 0
mem[72] = { 8'd48, 8'd10, 2'd1 }; // Age: 48, HR: 110, Class: 1
mem[73] = { 8'd57, 8'd44, 2'd2 }; // Age: 57, HR: 144, Class: 2
mem[74] = { 8'd44, 8'd79, 2'd0 }; // Age: 44, HR: 179, Class: 0
mem[75] = { 8'd45, 8'd47, 2'd3 }; // Age: 45, HR: 147, Class: 3
mem[76] = { 8'd45, 8'd48, 2'd0 }; // Age: 45, HR: 148, Class: 0
mem[77] = { 8'd49, 8'd40, 2'd1 }; // Age: 49, HR: 140, Class: 1
mem[78] = { 8'd46, 8'd20, 2'd0 }; // Age: 46, HR: 120, Class: 0
mem[79] = { 8'd67, 8'd8, 2'd2 }; // Age: 67, HR: 108, Class: 2
mem[80] = { 8'd47, 8'd45, 2'd0 }; // Age: 47, HR: 145, Class: 0
mem[81] = { 8'd52, 8'd24, 2'd1 }; // Age: 52, HR: 124, Class: 1
mem[82] = { 8'd54, 8'd56, 2'd0 }; // Age: 54, HR: 156, Class: 0
mem[83] = { 8'd69, 8'd18, 2'd2 }; // Age: 69, HR: 118, Class: 2
mem[84] = { 8'd62, 8'd242, 2'd0 }; // Age: 62, HR: 86, Class: 0
mem[85] = { 8'd58, 8'd50, 2'd0 }; // Age: 58, HR: 150, Class: 0
mem[86] = { 8'd64, 8'd14, 2'd1 }; // Age: 64, HR: 114, Class: 1
mem[87] = { 8'd48, 8'd18, 2'd0 }; // Age: 48, HR: 118, Class: 0
mem[88] = { 8'd59, 8'd17, 2'd1 }; // Age: 59, HR: 117, Class: 1
mem[89] = { 8'd44, 8'd50, 2'd1 }; // Age: 44, HR: 150, Class: 1
mem[90] = { 8'd77, 8'd62, 2'd3 }; // Age: 77, HR: 162, Class: 3
mem[91] = { 8'd64, 8'd54, 2'd0 }; // Age: 64, HR: 154, Class: 0
mem[92] = { 8'd42, 8'd50, 2'd0 }; // Age: 42, HR: 150, Class: 0
mem[93] = { 8'd54, 8'd54, 2'd1 }; // Age: 54, HR: 154, Class: 1
mem[94] = { 8'd70, 8'd29, 2'd2 }; // Age: 70, HR: 129, Class: 2
mem[95] = { 8'd61, 8'd38, 2'd1 }; // Age: 61, HR: 138, Class: 1
mem[96] = { 8'd54, 8'd37, 2'd0 }; // Age: 54, HR: 137, Class: 0
mem[97] = { 8'd55, 8'd37, 2'd0 }; // Age: 55, HR: 137, Class: 0
mem[98] = { 8'd60, 8'd41, 2'd3 }; // Age: 60, HR: 141, Class: 3
mem[99] = { 8'd58, 8'd5, 2'd1 }; // Age: 58, HR: 105, Class: 1
mem[100] = { 8'd64, 8'd45, 2'd1 }; // Age: 64, HR: 145, Class: 1
mem[101] = { 8'd41, 8'd82, 2'd0 }; // Age: 41, HR: 182, Class: 0
mem[102] = { 8'd65, 8'd5, 2'd3 }; // Age: 65, HR: 105, Class: 3
mem[103] = { 8'd44, 8'd27, 2'd0 }; // Age: 44, HR: 127, Class: 0
mem[104] = { 8'd64, 8'd22, 2'd3 }; // Age: 64, HR: 122, Class: 3
mem[105] = { 8'd39, 8'd20, 2'd0 }; // Age: 39, HR: 120, Class: 0
mem[106] = { 8'd44, 8'd53, 2'd2 }; // Age: 44, HR: 153, Class: 2
mem[107] = { 8'd40, 8'd236, 2'd0 }; // Age: 40, HR: 80, Class: 0
mem[108] = { 8'd46, 8'd72, 2'd0 }; // Age: 46, HR: 172, Class: 0
mem[109] = { 8'd53, 8'd6, 2'd1 }; // Age: 53, HR: 106, Class: 1
mem[110] = { 8'd66, 8'd20, 2'd2 }; // Age: 66, HR: 120, Class: 2
mem[111] = { 8'd45, 8'd40, 2'd0 }; // Age: 45, HR: 140, Class: 0
mem[112] = { 8'd34, 8'd80, 2'd1 }; // Age: 34, HR: 180, Class: 1
mem[113] = { 8'd65, 8'd14, 2'd3 }; // Age: 65, HR: 114, Class: 3
mem[114] = { 8'd51, 8'd73, 2'd1 }; // Age: 51, HR: 173, Class: 1
mem[115] = { 8'd52, 8'd62, 2'd0 }; // Age: 52, HR: 162, Class: 0
mem[116] = { 8'd57, 8'd0, 2'd0 }; // Age: 57, HR: 100, Class: 0
mem[117] = { 8'd54, 8'd13, 2'd2 }; // Age: 54, HR: 113, Class: 2
mem[118] = { 8'd68, 8'd51, 2'd0 }; // Age: 68, HR: 151, Class: 0
mem[119] = { 8'd69, 8'd240, 2'd2 }; // Age: 69, HR: 84, Class: 2
mem[120] = { 8'd55, 8'd30, 2'd1 }; // Age: 55, HR: 130, Class: 1
mem[121] = { 8'd40, 8'd50, 2'd0 }; // Age: 40, HR: 150, Class: 0
mem[122] = { 8'd44, 8'd70, 2'd0 }; // Age: 44, HR: 170, Class: 0
mem[123] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[124] = { 8'd56, 8'd28, 2'd0 }; // Age: 56, HR: 128, Class: 0
mem[125] = { 8'd58, 8'd31, 2'd1 }; // Age: 58, HR: 131, Class: 1
mem[126] = { 8'd35, 8'd30, 2'd1 }; // Age: 35, HR: 130, Class: 1
mem[127] = { 8'd38, 8'd34, 2'd1 }; // Age: 38, HR: 134, Class: 1
mem[128] = { 8'd54, 8'd0, 2'd1 }; // Age: 54, HR: 100, Class: 1
mem[129] = { 8'd47, 8'd74, 2'd0 }; // Age: 47, HR: 174, Class: 0
mem[130] = { 8'd60, 8'd10, 2'd3 }; // Age: 60, HR: 110, Class: 3
mem[131] = { 8'd51, 8'd70, 2'd0 }; // Age: 51, HR: 170, Class: 0
mem[132] = { 8'd56, 8'd63, 2'd0 }; // Age: 56, HR: 163, Class: 0
mem[133] = { 8'd45, 8'd10, 2'd0 }; // Age: 45, HR: 110, Class: 0
mem[134] = { 8'd67, 8'd25, 2'd3 }; // Age: 67, HR: 125, Class: 3
mem[135] = { 8'd62, 8'd52, 2'd0 }; // Age: 62, HR: 152, Class: 0
mem[136] = { 8'd52, 8'd69, 2'd0 }; // Age: 52, HR: 169, Class: 0
mem[137] = { 8'd65, 8'd14, 2'd3 }; // Age: 65, HR: 114, Class: 3
mem[138] = { 8'd66, 8'd14, 2'd0 }; // Age: 66, HR: 114, Class: 0
mem[139] = { 8'd43, 8'd65, 2'd0 }; // Age: 43, HR: 165, Class: 0
mem[140] = { 8'd50, 8'd59, 2'd0 }; // Age: 50, HR: 159, Class: 0
mem[141] = { 8'd57, 8'd20, 2'd1 }; // Age: 57, HR: 120, Class: 1
mem[142] = { 8'd49, 8'd45, 2'd2 }; // Age: 49, HR: 145, Class: 2
mem[143] = { 8'd64, 8'd58, 2'd1 }; // Age: 64, HR: 158, Class: 1
mem[144] = { 8'd50, 8'd28, 2'd3 }; // Age: 50, HR: 128, Class: 3
mem[145] = { 8'd43, 8'd30, 2'd1 }; // Age: 43, HR: 130, Class: 1
mem[146] = { 8'd49, 8'd35, 2'd0 }; // Age: 49, HR: 135, Class: 0
mem[147] = { 8'd56, 8'd50, 2'd1 }; // Age: 56, HR: 150, Class: 1
mem[148] = { 8'd60, 8'd57, 2'd1 }; // Age: 60, HR: 157, Class: 1
mem[149] = { 8'd50, 8'd20, 2'd1 }; // Age: 50, HR: 120, Class: 1
mem[150] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[151] = { 8'd61, 8'd15, 2'd3 }; // Age: 61, HR: 115, Class: 3
mem[152] = { 8'd60, 8'd40, 2'd0 }; // Age: 60, HR: 140, Class: 0
mem[153] = { 8'd54, 8'd18, 2'd1 }; // Age: 54, HR: 118, Class: 1
mem[154] = { 8'd64, 8'd6, 2'd1 }; // Age: 64, HR: 106, Class: 1
mem[155] = { 8'd43, 8'd40, 2'd2 }; // Age: 43, HR: 140, Class: 2
mem[156] = { 8'd55, 8'd37, 2'd0 }; // Age: 55, HR: 137, Class: 0
mem[157] = { 8'd53, 8'd35, 2'd2 }; // Age: 53, HR: 135, Class: 2
mem[158] = { 8'd57, 8'd48, 2'd1 }; // Age: 57, HR: 148, Class: 1
mem[159] = { 8'd41, 8'd72, 2'd0 }; // Age: 41, HR: 172, Class: 0
mem[160] = { 8'd46, 8'd52, 2'd0 }; // Age: 46, HR: 152, Class: 0
mem[161] = { 8'd43, 8'd30, 2'd1 }; // Age: 43, HR: 130, Class: 1
mem[162] = { 8'd59, 8'd20, 2'd1 }; // Age: 59, HR: 120, Class: 1
mem[163] = { 8'd48, 8'd10, 2'd0 }; // Age: 48, HR: 110, Class: 0
mem[164] = { 8'd63, 8'd244, 2'd3 }; // Age: 63, HR: 88, Class: 3
mem[165] = { 8'd47, 8'd25, 2'd0 }; // Age: 47, HR: 125, Class: 0
mem[166] = { 8'd58, 8'd30, 2'd3 }; // Age: 58, HR: 130, Class: 3
mem[167] = { 8'd52, 8'd62, 2'd0 }; // Age: 52, HR: 162, Class: 0
mem[168] = { 8'd51, 8'd252, 2'd0 }; // Age: 51, HR: 96, Class: 0
mem[169] = { 8'd41, 8'd30, 2'd1 }; // Age: 41, HR: 130, Class: 1
mem[170] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[171] = { 8'd62, 8'd34, 2'd1 }; // Age: 62, HR: 134, Class: 1
mem[172] = { 8'd56, 8'd24, 2'd1 }; // Age: 56, HR: 124, Class: 1
mem[173] = { 8'd55, 8'd0, 2'd2 }; // Age: 55, HR: 100, Class: 2
mem[174] = { 8'd60, 8'd40, 2'd1 }; // Age: 60, HR: 140, Class: 1
mem[175] = { 8'd41, 8'd53, 2'd0 }; // Age: 41, HR: 153, Class: 0
mem[176] = { 8'd52, 8'd252, 2'd1 }; // Age: 52, HR: 96, Class: 1
mem[177] = { 8'd52, 8'd61, 2'd1 }; // Age: 52, HR: 161, Class: 1
mem[178] = { 8'd63, 8'd240, 2'd3 }; // Age: 63, HR: 84, Class: 3
mem[179] = { 8'd59, 8'd40, 2'd0 }; // Age: 59, HR: 140, Class: 0
mem[180] = { 8'd49, 8'd35, 2'd0 }; // Age: 49, HR: 135, Class: 0
mem[181] = { 8'd52, 8'd69, 2'd0 }; // Age: 52, HR: 169, Class: 0
mem[182] = { 8'd64, 8'd22, 2'd3 }; // Age: 64, HR: 122, Class: 3
mem[183] = { 8'd56, 8'd238, 2'd1 }; // Age: 56, HR: 82, Class: 1
mem[184] = { 8'd70, 8'd12, 2'd3 }; // Age: 70, HR: 112, Class: 3
mem[185] = { 8'd52, 8'd50, 2'd1 }; // Age: 52, HR: 150, Class: 1
mem[186] = { 8'd42, 8'd78, 2'd0 }; // Age: 42, HR: 178, Class: 0
mem[187] = { 8'd60, 8'd25, 2'd1 }; // Age: 60, HR: 125, Class: 1
mem[188] = { 8'd68, 8'd51, 2'd0 }; // Age: 68, HR: 151, Class: 0
mem[189] = { 8'd69, 8'd240, 2'd2 }; // Age: 69, HR: 84, Class: 2
mem[190] = { 8'd63, 8'd54, 2'd3 }; // Age: 63, HR: 154, Class: 3
mem[191] = { 8'd49, 8'd63, 2'd0 }; // Age: 49, HR: 163, Class: 0
mem[192] = { 8'd44, 8'd80, 2'd0 }; // Age: 44, HR: 180, Class: 0
mem[193] = { 8'd62, 8'd50, 2'd1 }; // Age: 62, HR: 150, Class: 1
mem[194] = { 8'd59, 8'd25, 2'd1 }; // Age: 59, HR: 125, Class: 1
mem[195] = { 8'd61, 8'd13, 2'd1 }; // Age: 61, HR: 113, Class: 1
mem[196] = { 8'd44, 8'd0, 2'd1 }; // Age: 44, HR: 100, Class: 1
mem[197] = { 8'd56, 8'd50, 2'd1 }; // Age: 56, HR: 150, Class: 1
mem[198] = { 8'd54, 8'd10, 2'd3 }; // Age: 54, HR: 110, Class: 3
mem[199] = { 8'd62, 8'd50, 2'd1 }; // Age: 62, HR: 150, Class: 1
mem[200] = { 8'd66, 8'd14, 2'd0 }; // Age: 66, HR: 114, Class: 0
mem[201] = { 8'd47, 8'd24, 2'd1 }; // Age: 47, HR: 124, Class: 1
mem[202] = { 8'd44, 8'd50, 2'd1 }; // Age: 44, HR: 150, Class: 1
mem[203] = { 8'd39, 8'd70, 2'd0 }; // Age: 39, HR: 170, Class: 0
mem[204] = { 8'd63, 8'd60, 2'd0 }; // Age: 63, HR: 160, Class: 0
mem[205] = { 8'd38, 8'd29, 2'd0 }; // Age: 38, HR: 129, Class: 0
mem[206] = { 8'd53, 8'd22, 2'd1 }; // Age: 53, HR: 122, Class: 1
mem[207] = { 8'd46, 8'd25, 2'd1 }; // Age: 46, HR: 125, Class: 1
mem[208] = { 8'd40, 8'd88, 2'd0 }; // Age: 40, HR: 188, Class: 0
mem[209] = { 8'd56, 8'd40, 2'd0 }; // Age: 56, HR: 140, Class: 0
mem[210] = { 8'd52, 8'd69, 2'd0 }; // Age: 52, HR: 169, Class: 0
mem[211] = { 8'd69, 8'd46, 2'd2 }; // Age: 69, HR: 146, Class: 2
mem[212] = { 8'd63, 8'd69, 2'd1 }; // Age: 63, HR: 169, Class: 1
mem[213] = { 8'd46, 8'd16, 2'd0 }; // Age: 46, HR: 116, Class: 0
mem[214] = { 8'd45, 8'd44, 2'd0 }; // Age: 45, HR: 144, Class: 0
mem[215] = { 8'd55, 8'd30, 2'd3 }; // Age: 55, HR: 130, Class: 3
mem[216] = { 8'd52, 8'd20, 2'd2 }; // Age: 52, HR: 120, Class: 2
mem[217] = { 8'd51, 8'd4, 2'd3 }; // Age: 51, HR: 104, Class: 3
mem[218] = { 8'd77, 8'd10, 2'd3 }; // Age: 77, HR: 110, Class: 3
mem[219] = { 8'd70, 8'd43, 2'd0 }; // Age: 70, HR: 143, Class: 0
mem[220] = { 8'd42, 8'd36, 2'd0 }; // Age: 42, HR: 136, Class: 0
mem[221] = { 8'd67, 8'd25, 2'd2 }; // Age: 67, HR: 125, Class: 2
mem[222] = { 8'd54, 8'd37, 2'd0 }; // Age: 54, HR: 137, Class: 0
mem[223] = { 8'd49, 8'd30, 2'd0 }; // Age: 49, HR: 130, Class: 0
mem[224] = { 8'd55, 8'd55, 2'd1 }; // Age: 55, HR: 155, Class: 1
mem[225] = { 8'd35, 8'd80, 2'd0 }; // Age: 35, HR: 180, Class: 0
mem[226] = { 8'd60, 8'd219, 2'd3 }; // Age: 60, HR: 63, Class: 3
mem[227] = { 8'd63, 8'd69, 2'd1 }; // Age: 63, HR: 169, Class: 1
mem[228] = { 8'd61, 8'd0, 2'd3 }; // Age: 61, HR: 100, Class: 3
mem[229] = { 8'd74, 8'd21, 2'd0 }; // Age: 74, HR: 121, Class: 0
mem[230] = { 8'd61, 8'd15, 2'd3 }; // Age: 61, HR: 115, Class: 3
mem[231] = { 8'd57, 8'd254, 2'd2 }; // Age: 57, HR: 98, Class: 2
mem[232] = { 8'd59, 8'd54, 2'd0 }; // Age: 59, HR: 154, Class: 0
mem[233] = { 8'd44, 8'd70, 2'd0 }; // Age: 44, HR: 170, Class: 0
mem[234] = { 8'd59, 8'd19, 2'd1 }; // Age: 59, HR: 119, Class: 1
mem[235] = { 8'd41, 8'd76, 2'd2 }; // Age: 41, HR: 176, Class: 2
mem[236] = { 8'd56, 8'd28, 2'd0 }; // Age: 56, HR: 128, Class: 0
mem[237] = { 8'd49, 8'd26, 2'd1 }; // Age: 49, HR: 126, Class: 1
mem[238] = { 8'd62, 8'd228, 2'd3 }; // Age: 62, HR: 72, Class: 3
mem[239] = { 8'd52, 8'd90, 2'd0 }; // Age: 52, HR: 190, Class: 0
mem[240] = { 8'd71, 8'd15, 2'd3 }; // Age: 71, HR: 115, Class: 3
mem[241] = { 8'd38, 8'd66, 2'd1 }; // Age: 38, HR: 166, Class: 1
mem[242] = { 8'd53, 8'd55, 2'd0 }; // Age: 53, HR: 155, Class: 0
mem[243] = { 8'd52, 8'd252, 2'd1 }; // Age: 52, HR: 96, Class: 1
mem[244] = { 8'd59, 8'd34, 2'd2 }; // Age: 59, HR: 134, Class: 2
mem[245] = { 8'd48, 8'd15, 2'd1 }; // Age: 48, HR: 115, Class: 1
mem[246] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[247] = { 8'd46, 8'd40, 2'd0 }; // Age: 46, HR: 140, Class: 0
mem[248] = { 8'd46, 8'd40, 2'd0 }; // Age: 46, HR: 140, Class: 0
mem[249] = { 8'd52, 8'd90, 2'd0 }; // Age: 52, HR: 190, Class: 0
mem[250] = { 8'd43, 8'd40, 2'd2 }; // Age: 43, HR: 140, Class: 2
mem[251] = { 8'd50, 8'd39, 2'd1 }; // Age: 50, HR: 139, Class: 1
mem[252] = { 8'd45, 8'd48, 2'd0 }; // Age: 45, HR: 148, Class: 0
mem[253] = { 8'd63, 8'd54, 2'd3 }; // Age: 63, HR: 154, Class: 3
mem[254] = { 8'd52, 8'd90, 2'd0 }; // Age: 52, HR: 190, Class: 0
mem[255] = { 8'd67, 8'd8, 2'd2 }; // Age: 67, HR: 108, Class: 2
mem[256] = { 8'd53, 8'd20, 2'd3 }; // Age: 53, HR: 120, Class: 3
mem[257] = { 8'd59, 8'd82, 2'd0 }; // Age: 59, HR: 182, Class: 0
mem[258] = { 8'd52, 8'd24, 2'd1 }; // Age: 52, HR: 124, Class: 1
mem[259] = { 8'd58, 8'd18, 2'd2 }; // Age: 58, HR: 118, Class: 2
mem[260] = { 8'd63, 8'd20, 2'd0 }; // Age: 63, HR: 120, Class: 0
mem[261] = { 8'd63, 8'd69, 2'd1 }; // Age: 63, HR: 169, Class: 1
mem[262] = { 8'd46, 8'd16, 2'd0 }; // Age: 46, HR: 116, Class: 0
mem[263] = { 8'd48, 8'd38, 2'd0 }; // Age: 48, HR: 138, Class: 0
mem[264] = { 8'd53, 8'd20, 2'd0 }; // Age: 53, HR: 120, Class: 0
mem[265] = { 8'd62, 8'd63, 2'd0 }; // Age: 62, HR: 163, Class: 0
mem[266] = { 8'd44, 8'd53, 2'd2 }; // Age: 44, HR: 153, Class: 2
mem[267] = { 8'd61, 8'd15, 2'd3 }; // Age: 61, HR: 115, Class: 3
mem[268] = { 8'd59, 8'd17, 2'd1 }; // Age: 59, HR: 117, Class: 1
mem[269] = { 8'd59, 8'd19, 2'd1 }; // Age: 59, HR: 119, Class: 1
mem[270] = { 8'd67, 8'd25, 2'd2 }; // Age: 67, HR: 125, Class: 2
mem[271] = { 8'd50, 8'd16, 2'd0 }; // Age: 50, HR: 116, Class: 0
mem[272] = { 8'd58, 8'd56, 2'd2 }; // Age: 58, HR: 156, Class: 2
mem[273] = { 8'd62, 8'd20, 2'd3 }; // Age: 62, HR: 120, Class: 3
mem[274] = { 8'd53, 8'd40, 2'd0 }; // Age: 53, HR: 140, Class: 0
mem[275] = { 8'd57, 8'd73, 2'd0 }; // Age: 57, HR: 173, Class: 0
mem[276] = { 8'd59, 8'd45, 2'd0 }; // Age: 59, HR: 145, Class: 0
mem[277] = { 8'd51, 8'd43, 2'd0 }; // Age: 51, HR: 143, Class: 0
mem[278] = { 8'd48, 8'd60, 2'd0 }; // Age: 48, HR: 160, Class: 0
mem[279] = { 8'd59, 8'd20, 2'd1 }; // Age: 59, HR: 120, Class: 1
mem[280] = { 8'd63, 8'd44, 2'd2 }; // Age: 63, HR: 144, Class: 2
mem[281] = { 8'd58, 8'd31, 2'd0 }; // Age: 58, HR: 131, Class: 0
mem[282] = { 8'd57, 8'd19, 2'd3 }; // Age: 57, HR: 119, Class: 3
mem[283] = { 8'd42, 8'd255, 2'd2 }; // Age: 42, HR: 99, Class: 2
mem[284] = { 8'd45, 8'd52, 2'd0 }; // Age: 45, HR: 152, Class: 0
mem[285] = { 8'd48, 8'd3, 2'd1 }; // Age: 48, HR: 103, Class: 1
mem[286] = { 8'd61, 8'd236, 2'd3 }; // Age: 61, HR: 80, Class: 3
mem[287] = { 8'd64, 8'd31, 2'd1 }; // Age: 64, HR: 131, Class: 1
mem[288] = { 8'd42, 8'd28, 2'd1 }; // Age: 42, HR: 128, Class: 1
mem[289] = { 8'd50, 8'd59, 2'd0 }; // Age: 50, HR: 159, Class: 0
mem[290] = { 8'd55, 8'd11, 2'd3 }; // Age: 55, HR: 111, Class: 3
mem[291] = { 8'd42, 8'd94, 2'd0 }; // Age: 42, HR: 194, Class: 0
mem[292] = { 8'd37, 8'd84, 2'd0 }; // Age: 37, HR: 184, Class: 0
mem[293] = { 8'd55, 8'd55, 2'd0 }; // Age: 55, HR: 155, Class: 0
mem[294] = { 8'd41, 8'd42, 2'd0 }; // Age: 41, HR: 142, Class: 0
mem[295] = { 8'd58, 8'd10, 2'd2 }; // Age: 58, HR: 110, Class: 2
mem[296] = { 8'd57, 8'd48, 2'd1 }; // Age: 57, HR: 148, Class: 1
mem[297] = { 8'd53, 8'd6, 2'd1 }; // Age: 53, HR: 106, Class: 1
mem[298] = { 8'd48, 8'd38, 2'd0 }; // Age: 48, HR: 138, Class: 0
mem[299] = { 8'd40, 8'd38, 2'd0 }; // Age: 40, HR: 138, Class: 0
mem[300] = { 8'd48, 8'd3, 2'd1 }; // Age: 48, HR: 103, Class: 1
mem[301] = { 8'd57, 8'd24, 2'd3 }; // Age: 57, HR: 124, Class: 3
mem[302] = { 8'd41, 8'd79, 2'd0 }; // Age: 41, HR: 179, Class: 0
mem[303] = { 8'd55, 8'd0, 2'd2 }; // Age: 55, HR: 100, Class: 2
mem[304] = { 8'd68, 8'd20, 2'd3 }; // Age: 68, HR: 120, Class: 3
mem[305] = { 8'd66, 8'd40, 2'd1 }; // Age: 66, HR: 140, Class: 1
mem[306] = { 8'd62, 8'd16, 2'd0 }; // Age: 62, HR: 116, Class: 0
mem[307] = { 8'd53, 8'd22, 2'd1 }; // Age: 53, HR: 122, Class: 1
mem[308] = { 8'd57, 8'd248, 2'd1 }; // Age: 57, HR: 92, Class: 1
mem[309] = { 8'd39, 8'd20, 2'd0 }; // Age: 39, HR: 120, Class: 0
mem[310] = { 8'd53, 8'd20, 2'd1 }; // Age: 53, HR: 120, Class: 1
mem[311] = { 8'd75, 8'd8, 2'd1 }; // Age: 75, HR: 108, Class: 1
mem[312] = { 8'd56, 8'd40, 2'd0 }; // Age: 56, HR: 140, Class: 0
mem[313] = { 8'd52, 8'd78, 2'd0 }; // Age: 52, HR: 178, Class: 0
mem[314] = { 8'd50, 8'd70, 2'd0 }; // Age: 50, HR: 170, Class: 0
mem[315] = { 8'd57, 8'd23, 2'd1 }; // Age: 57, HR: 123, Class: 1
mem[316] = { 8'd43, 8'd22, 2'd3 }; // Age: 43, HR: 122, Class: 3
mem[317] = { 8'd60, 8'd71, 2'd0 }; // Age: 60, HR: 171, Class: 0
mem[318] = { 8'd53, 8'd6, 2'd1 }; // Age: 53, HR: 106, Class: 1
mem[319] = { 8'd64, 8'd31, 2'd1 }; // Age: 64, HR: 131, Class: 1
mem[320] = { 8'd40, 8'd38, 2'd0 }; // Age: 40, HR: 138, Class: 0
mem[321] = { 8'd50, 8'd56, 2'd3 }; // Age: 50, HR: 156, Class: 3
mem[322] = { 8'd55, 8'd43, 2'd1 }; // Age: 55, HR: 143, Class: 1
mem[323] = { 8'd67, 8'd8, 2'd2 }; // Age: 67, HR: 108, Class: 2
mem[324] = { 8'd28, 8'd85, 2'd0 }; // Age: 28, HR: 185, Class: 0
mem[325] = { 8'd51, 8'd57, 2'd0 }; // Age: 51, HR: 157, Class: 0
mem[326] = { 8'd56, 8'd253, 2'd0 }; // Age: 56, HR: 97, Class: 0
mem[327] = { 8'd54, 8'd10, 2'd0 }; // Age: 54, HR: 110, Class: 0
mem[328] = { 8'd43, 8'd20, 2'd3 }; // Age: 43, HR: 120, Class: 3
mem[329] = { 8'd68, 8'd51, 2'd0 }; // Age: 68, HR: 151, Class: 0
mem[330] = { 8'd63, 8'd47, 2'd2 }; // Age: 63, HR: 147, Class: 2
mem[331] = { 8'd49, 8'd26, 2'd1 }; // Age: 49, HR: 126, Class: 1
mem[332] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[333] = { 8'd56, 8'd21, 2'd1 }; // Age: 56, HR: 121, Class: 1
mem[334] = { 8'd70, 8'd29, 2'd2 }; // Age: 70, HR: 129, Class: 2
mem[335] = { 8'd50, 8'd26, 2'd3 }; // Age: 50, HR: 126, Class: 3
mem[336] = { 8'd54, 8'd47, 2'd0 }; // Age: 54, HR: 147, Class: 0
mem[337] = { 8'd49, 8'd60, 2'd0 }; // Age: 49, HR: 160, Class: 0
mem[338] = { 8'd42, 8'd22, 2'd0 }; // Age: 42, HR: 122, Class: 0
mem[339] = { 8'd44, 8'd88, 2'd0 }; // Age: 44, HR: 188, Class: 0
mem[340] = { 8'd65, 8'd27, 2'd2 }; // Age: 65, HR: 127, Class: 2
mem[341] = { 8'd59, 8'd15, 2'd1 }; // Age: 59, HR: 115, Class: 1
mem[342] = { 8'd51, 8'd4, 2'd3 }; // Age: 51, HR: 104, Class: 3
mem[343] = { 8'd49, 8'd252, 2'd1 }; // Age: 49, HR: 96, Class: 1
mem[344] = { 8'd50, 8'd39, 2'd1 }; // Age: 50, HR: 139, Class: 1
mem[345] = { 8'd51, 8'd20, 2'd0 }; // Age: 51, HR: 120, Class: 0
mem[346] = { 8'd51, 8'd20, 2'd0 }; // Age: 51, HR: 120, Class: 0
mem[347] = { 8'd71, 8'd30, 2'd0 }; // Age: 71, HR: 130, Class: 0
mem[348] = { 8'd56, 8'd254, 2'd1 }; // Age: 56, HR: 98, Class: 1
mem[349] = { 8'd51, 8'd57, 2'd0 }; // Age: 51, HR: 157, Class: 0
mem[350] = { 8'd47, 8'd43, 2'd0 }; // Age: 47, HR: 143, Class: 0
mem[351] = { 8'd56, 8'd44, 2'd1 }; // Age: 56, HR: 144, Class: 1
mem[352] = { 8'd48, 8'd15, 2'd1 }; // Age: 48, HR: 115, Class: 1
mem[353] = { 8'd56, 8'd40, 2'd0 }; // Age: 56, HR: 140, Class: 0
mem[354] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[355] = { 8'd67, 8'd60, 2'd0 }; // Age: 67, HR: 160, Class: 0
mem[356] = { 8'd62, 8'd38, 2'd1 }; // Age: 62, HR: 138, Class: 1
mem[357] = { 8'd39, 8'd20, 2'd0 }; // Age: 39, HR: 120, Class: 0
mem[358] = { 8'd65, 8'd54, 2'd0 }; // Age: 65, HR: 154, Class: 0
mem[359] = { 8'd62, 8'd242, 2'd0 }; // Age: 62, HR: 86, Class: 0
mem[360] = { 8'd54, 8'd58, 2'd0 }; // Age: 54, HR: 158, Class: 0
mem[361] = { 8'd44, 8'd27, 2'd0 }; // Age: 44, HR: 127, Class: 0
mem[362] = { 8'd61, 8'd10, 2'd1 }; // Age: 61, HR: 110, Class: 1
mem[363] = { 8'd46, 8'd56, 2'd0 }; // Age: 46, HR: 156, Class: 0
mem[364] = { 8'd65, 8'd12, 2'd1 }; // Age: 65, HR: 112, Class: 1
mem[365] = { 8'd48, 8'd10, 2'd1 }; // Age: 48, HR: 110, Class: 1
mem[366] = { 8'd48, 8'd10, 2'd0 }; // Age: 48, HR: 110, Class: 0
mem[367] = { 8'd66, 8'd52, 2'd0 }; // Age: 66, HR: 152, Class: 0
mem[368] = { 8'd70, 8'd29, 2'd2 }; // Age: 70, HR: 129, Class: 2
mem[369] = { 8'd46, 8'd50, 2'd1 }; // Age: 46, HR: 150, Class: 1
mem[370] = { 8'd47, 8'd74, 2'd0 }; // Age: 47, HR: 174, Class: 0
mem[371] = { 8'd43, 8'd65, 2'd0 }; // Age: 43, HR: 165, Class: 0
mem[372] = { 8'd68, 8'd15, 2'd0 }; // Age: 68, HR: 115, Class: 0
mem[373] = { 8'd48, 8'd60, 2'd0 }; // Age: 48, HR: 160, Class: 0
mem[374] = { 8'd53, 8'd22, 2'd1 }; // Age: 53, HR: 122, Class: 1
mem[375] = { 8'd64, 8'd58, 2'd1 }; // Age: 64, HR: 158, Class: 1
mem[376] = { 8'd61, 8'd45, 2'd2 }; // Age: 61, HR: 145, Class: 2
mem[377] = { 8'd55, 8'd55, 2'd0 }; // Age: 55, HR: 155, Class: 0
mem[378] = { 8'd56, 8'd0, 2'd0 }; // Age: 56, HR: 100, Class: 0
mem[379] = { 8'd45, 8'd70, 2'd0 }; // Age: 45, HR: 170, Class: 0
mem[380] = { 8'd58, 8'd62, 2'd0 }; // Age: 58, HR: 162, Class: 0
mem[381] = { 8'd60, 8'd33, 2'd0 }; // Age: 60, HR: 133, Class: 0
mem[382] = { 8'd59, 8'd250, 2'd3 }; // Age: 59, HR: 94, Class: 3
mem[383] = { 8'd57, 8'd12, 2'd1 }; // Age: 57, HR: 112, Class: 1
mem[384] = { 8'd66, 8'd32, 2'd2 }; // Age: 66, HR: 132, Class: 2
mem[385] = { 8'd43, 8'd75, 2'd0 }; // Age: 43, HR: 175, Class: 0
mem[386] = { 8'd51, 8'd50, 2'd1 }; // Age: 51, HR: 150, Class: 1
mem[387] = { 8'd53, 8'd62, 2'd0 }; // Age: 53, HR: 162, Class: 0
mem[388] = { 8'd57, 8'd44, 2'd2 }; // Age: 57, HR: 144, Class: 2
mem[389] = { 8'd55, 8'd30, 2'd3 }; // Age: 55, HR: 130, Class: 3
mem[390] = { 8'd58, 8'd72, 2'd0 }; // Age: 58, HR: 172, Class: 0
mem[391] = { 8'd34, 8'd92, 2'd0 }; // Age: 34, HR: 192, Class: 0
mem[392] = { 8'd66, 8'd52, 2'd0 }; // Age: 66, HR: 152, Class: 0
mem[393] = { 8'd63, 8'd60, 2'd0 }; // Age: 63, HR: 160, Class: 0
mem[394] = { 8'd42, 8'd28, 2'd1 }; // Age: 42, HR: 128, Class: 1
mem[395] = { 8'd35, 8'd74, 2'd0 }; // Age: 35, HR: 174, Class: 0
mem[396] = { 8'd59, 8'd24, 2'd0 }; // Age: 59, HR: 124, Class: 0
mem[397] = { 8'd54, 8'd10, 2'd0 }; // Age: 54, HR: 110, Class: 0
mem[398] = { 8'd41, 8'd28, 2'd0 }; // Age: 41, HR: 128, Class: 0
mem[399] = { 8'd70, 8'd29, 2'd2 }; // Age: 70, HR: 129, Class: 2
mem[400] = { 8'd56, 8'd21, 2'd1 }; // Age: 56, HR: 121, Class: 1
mem[401] = { 8'd50, 8'd50, 2'd1 }; // Age: 50, HR: 150, Class: 1
mem[402] = { 8'd54, 8'd18, 2'd1 }; // Age: 54, HR: 118, Class: 1
mem[403] = { 8'd51, 8'd22, 2'd3 }; // Age: 51, HR: 122, Class: 3
mem[404] = { 8'd65, 8'd57, 2'd0 }; // Age: 65, HR: 157, Class: 0
mem[405] = { 8'd49, 8'd56, 2'd1 }; // Age: 49, HR: 156, Class: 1
mem[406] = { 8'd48, 8'd68, 2'd1 }; // Age: 48, HR: 168, Class: 1
mem[407] = { 8'd53, 8'd11, 2'd0 }; // Age: 53, HR: 111, Class: 0
mem[408] = { 8'd59, 8'd82, 2'd0 }; // Age: 59, HR: 182, Class: 0
mem[409] = { 8'd58, 8'd71, 2'd1 }; // Age: 58, HR: 171, Class: 1
mem[410] = { 8'd58, 8'd50, 2'd0 }; // Age: 58, HR: 150, Class: 0
mem[411] = { 8'd58, 8'd65, 2'd3 }; // Age: 58, HR: 165, Class: 3
mem[412] = { 8'd44, 8'd35, 2'd0 }; // Age: 44, HR: 135, Class: 0
mem[413] = { 8'd52, 8'd20, 2'd1 }; // Age: 52, HR: 120, Class: 1
mem[414] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[415] = { 8'd77, 8'd10, 2'd3 }; // Age: 77, HR: 110, Class: 3
mem[416] = { 8'd43, 8'd20, 2'd3 }; // Age: 43, HR: 120, Class: 3
mem[417] = { 8'd58, 8'd31, 2'd0 }; // Age: 58, HR: 131, Class: 0
mem[418] = { 8'd41, 8'd42, 2'd0 }; // Age: 41, HR: 142, Class: 0
mem[419] = { 8'd38, 8'd66, 2'd1 }; // Age: 38, HR: 166, Class: 1
mem[420] = { 8'd57, 8'd74, 2'd1 }; // Age: 57, HR: 174, Class: 1
mem[421] = { 8'd48, 8'd66, 2'd3 }; // Age: 48, HR: 166, Class: 3
mem[422] = { 8'd40, 8'd44, 2'd2 }; // Age: 40, HR: 144, Class: 2
mem[423] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[424] = { 8'd63, 8'd254, 2'd1 }; // Age: 63, HR: 98, Class: 1
mem[425] = { 8'd41, 8'd32, 2'd0 }; // Age: 41, HR: 132, Class: 0
mem[426] = { 8'd50, 8'd63, 2'd0 }; // Age: 50, HR: 163, Class: 0
mem[427] = { 8'd64, 8'd5, 2'd0 }; // Age: 64, HR: 105, Class: 0
mem[428] = { 8'd46, 8'd56, 2'd0 }; // Age: 46, HR: 156, Class: 0
mem[429] = { 8'd42, 8'd73, 2'd0 }; // Age: 42, HR: 173, Class: 0
mem[430] = { 8'd36, 8'd72, 2'd0 }; // Age: 36, HR: 172, Class: 0
mem[431] = { 8'd54, 8'd26, 2'd3 }; // Age: 54, HR: 126, Class: 3
mem[432] = { 8'd54, 8'd60, 2'd0 }; // Age: 54, HR: 160, Class: 0
mem[433] = { 8'd67, 8'd50, 2'd3 }; // Age: 67, HR: 150, Class: 3
mem[434] = { 8'd46, 8'd25, 2'd1 }; // Age: 46, HR: 125, Class: 1
mem[435] = { 8'd52, 8'd24, 2'd1 }; // Age: 52, HR: 124, Class: 1
mem[436] = { 8'd54, 8'd5, 2'd1 }; // Age: 54, HR: 105, Class: 1
mem[437] = { 8'd36, 8'd72, 2'd0 }; // Age: 36, HR: 172, Class: 0
mem[438] = { 8'd61, 8'd5, 2'd1 }; // Age: 61, HR: 105, Class: 1
mem[439] = { 8'd40, 8'd236, 2'd0 }; // Age: 40, HR: 80, Class: 0
mem[440] = { 8'd51, 8'd27, 2'd2 }; // Age: 51, HR: 127, Class: 2
mem[441] = { 8'd58, 8'd44, 2'd0 }; // Age: 58, HR: 144, Class: 0
mem[442] = { 8'd61, 8'd254, 2'd3 }; // Age: 61, HR: 98, Class: 3
mem[443] = { 8'd57, 8'd0, 2'd3 }; // Age: 57, HR: 100, Class: 3
mem[444] = { 8'd53, 8'd15, 2'd1 }; // Age: 53, HR: 115, Class: 1
mem[445] = { 8'd64, 8'd252, 2'd3 }; // Age: 64, HR: 96, Class: 3
mem[446] = { 8'd62, 8'd52, 2'd0 }; // Age: 62, HR: 152, Class: 0
mem[447] = { 8'd46, 8'd40, 2'd0 }; // Age: 46, HR: 140, Class: 0
mem[448] = { 8'd67, 8'd30, 2'd2 }; // Age: 67, HR: 130, Class: 2
mem[449] = { 8'd71, 8'd30, 2'd0 }; // Age: 71, HR: 130, Class: 0
mem[450] = { 8'd47, 8'd25, 2'd0 }; // Age: 47, HR: 125, Class: 0
mem[451] = { 8'd74, 8'd30, 2'd3 }; // Age: 74, HR: 130, Class: 3
mem[452] = { 8'd67, 8'd227, 2'd2 }; // Age: 67, HR: 71, Class: 2
mem[453] = { 8'd57, 8'd244, 2'd1 }; // Age: 57, HR: 88, Class: 1
mem[454] = { 8'd55, 8'd32, 2'd3 }; // Age: 55, HR: 132, Class: 3
mem[455] = { 8'd58, 8'd50, 2'd0 }; // Age: 58, HR: 150, Class: 0
mem[456] = { 8'd61, 8'd13, 2'd1 }; // Age: 61, HR: 113, Class: 1
mem[457] = { 8'd59, 8'd28, 2'd2 }; // Age: 59, HR: 128, Class: 2
mem[458] = { 8'd48, 8'd248, 2'd1 }; // Age: 48, HR: 92, Class: 1
mem[459] = { 8'd48, 8'd62, 2'd1 }; // Age: 48, HR: 162, Class: 1
mem[460] = { 8'd49, 8'd74, 2'd0 }; // Age: 49, HR: 174, Class: 0
mem[461] = { 8'd60, 8'd25, 2'd1 }; // Age: 60, HR: 125, Class: 1
mem[462] = { 8'd57, 8'd60, 2'd3 }; // Age: 57, HR: 160, Class: 3
mem[463] = { 8'd46, 8'd25, 2'd1 }; // Age: 46, HR: 125, Class: 1
mem[464] = { 8'd75, 8'd12, 2'd0 }; // Age: 75, HR: 112, Class: 0
mem[465] = { 8'd42, 8'd78, 2'd0 }; // Age: 42, HR: 178, Class: 0
mem[466] = { 8'd61, 8'd233, 2'd3 }; // Age: 61, HR: 77, Class: 3
mem[467] = { 8'd49, 8'd71, 2'd0 }; // Age: 49, HR: 171, Class: 0
mem[468] = { 8'd36, 8'd84, 2'd0 }; // Age: 36, HR: 184, Class: 0
mem[469] = { 8'd57, 8'd44, 2'd2 }; // Age: 57, HR: 144, Class: 2
mem[470] = { 8'd49, 8'd56, 2'd1 }; // Age: 49, HR: 156, Class: 1
mem[471] = { 8'd48, 8'd0, 2'd0 }; // Age: 48, HR: 100, Class: 0
mem[472] = { 8'd56, 8'd255, 2'd2 }; // Age: 56, HR: 99, Class: 2
mem[473] = { 8'd56, 8'd14, 2'd0 }; // Age: 56, HR: 114, Class: 0
mem[474] = { 8'd52, 8'd84, 2'd0 }; // Age: 52, HR: 184, Class: 0
mem[475] = { 8'd62, 8'd45, 2'd3 }; // Age: 62, HR: 145, Class: 3
mem[476] = { 8'd41, 8'd44, 2'd0 }; // Age: 41, HR: 144, Class: 0
mem[477] = { 8'd64, 8'd35, 2'd2 }; // Age: 64, HR: 135, Class: 2
mem[478] = { 8'd65, 8'd20, 2'd3 }; // Age: 65, HR: 120, Class: 3
mem[479] = { 8'd60, 8'd41, 2'd3 }; // Age: 60, HR: 141, Class: 3
mem[480] = { 8'd61, 8'd254, 2'd3 }; // Age: 61, HR: 98, Class: 3
mem[481] = { 8'd41, 8'd68, 2'd0 }; // Age: 41, HR: 168, Class: 0
mem[482] = { 8'd57, 8'd82, 2'd1 }; // Age: 57, HR: 182, Class: 1
mem[483] = { 8'd63, 8'd242, 2'd3 }; // Age: 63, HR: 86, Class: 3
mem[484] = { 8'd56, 8'd24, 2'd1 }; // Age: 56, HR: 124, Class: 1
mem[485] = { 8'd69, 8'd46, 2'd2 }; // Age: 69, HR: 146, Class: 2
mem[486] = { 8'd65, 8'd74, 2'd1 }; // Age: 65, HR: 174, Class: 1
mem[487] = { 8'd60, 8'd60, 2'd0 }; // Age: 60, HR: 160, Class: 0
mem[488] = { 8'd34, 8'd68, 2'd0 }; // Age: 34, HR: 168, Class: 0
mem[489] = { 8'd54, 8'd5, 2'd1 }; // Age: 54, HR: 105, Class: 1
mem[490] = { 8'd39, 8'd32, 2'd0 }; // Age: 39, HR: 132, Class: 0
mem[491] = { 8'd29, 8'd60, 2'd0 }; // Age: 29, HR: 160, Class: 0
mem[492] = { 8'd62, 8'd228, 2'd3 }; // Age: 62, HR: 72, Class: 3
mem[493] = { 8'd61, 8'd13, 2'd1 }; // Age: 61, HR: 113, Class: 1
mem[494] = { 8'd48, 8'd59, 2'd3 }; // Age: 48, HR: 159, Class: 3
mem[495] = { 8'd58, 8'd225, 2'd0 }; // Age: 58, HR: 69, Class: 0
mem[496] = { 8'd44, 8'd88, 2'd0 }; // Age: 44, HR: 188, Class: 0
mem[497] = { 8'd54, 8'd40, 2'd0 }; // Age: 54, HR: 140, Class: 0
mem[498] = { 8'd43, 8'd40, 2'd2 }; // Age: 43, HR: 140, Class: 2
mem[499] = { 8'd44, 8'd69, 2'd0 }; // Age: 44, HR: 169, Class: 0
mem[500] = { 8'd44, 8'd53, 2'd2 }; // Age: 44, HR: 153, Class: 2
mem[501] = { 8'd55, 8'd43, 2'd1 }; // Age: 55, HR: 143, Class: 1
mem[502] = { 8'd47, 8'd24, 2'd1 }; // Age: 47, HR: 124, Class: 1
mem[503] = { 8'd41, 8'd72, 2'd0 }; // Age: 41, HR: 172, Class: 0
mem[504] = { 8'd57, 8'd59, 2'd0 }; // Age: 57, HR: 159, Class: 0
mem[505] = { 8'd67, 8'd25, 2'd3 }; // Age: 67, HR: 125, Class: 3
mem[506] = { 8'd58, 8'd6, 2'd1 }; // Age: 58, HR: 106, Class: 1
mem[507] = { 8'd41, 8'd80, 2'd0 }; // Age: 41, HR: 180, Class: 0
mem[508] = { 8'd51, 8'd23, 2'd0 }; // Age: 51, HR: 123, Class: 0
mem[509] = { 8'd53, 8'd60, 2'd0 }; // Age: 53, HR: 160, Class: 0
mem[510] = { 8'd66, 8'd40, 2'd1 }; // Age: 66, HR: 140, Class: 1
mem[511] = { 8'd56, 8'd0, 2'd2 }; // Age: 56, HR: 100, Class: 2
mem[512] = { 8'd40, 8'd81, 2'd1 }; // Age: 40, HR: 181, Class: 1
mem[513] = { 8'd43, 8'd38, 2'd0 }; // Age: 43, HR: 138, Class: 0
mem[514] = { 8'd52, 8'd238, 2'd2 }; // Age: 52, HR: 82, Class: 2
mem[515] = { 8'd54, 8'd56, 2'd0 }; // Age: 54, HR: 156, Class: 0
mem[516] = { 8'd59, 8'd250, 2'd3 }; // Age: 59, HR: 94, Class: 3
mem[517] = { 8'd56, 8'd21, 2'd1 }; // Age: 56, HR: 121, Class: 1
mem[518] = { 8'd56, 8'd48, 2'd2 }; // Age: 56, HR: 148, Class: 2
mem[519] = { 8'd65, 8'd27, 2'd2 }; // Age: 65, HR: 127, Class: 2
mem[520] = { 8'd38, 8'd5, 2'd1 }; // Age: 38, HR: 105, Class: 1
mem[521] = { 8'd65, 8'd40, 2'd3 }; // Age: 65, HR: 140, Class: 3
mem[522] = { 8'd38, 8'd28, 2'd1 }; // Age: 38, HR: 128, Class: 1
mem[523] = { 8'd41, 8'd58, 2'd1 }; // Age: 41, HR: 158, Class: 1
mem[524] = { 8'd40, 8'd38, 2'd0 }; // Age: 40, HR: 138, Class: 0
mem[525] = { 8'd52, 8'd80, 2'd2 }; // Age: 52, HR: 180, Class: 2
mem[526] = { 8'd57, 8'd254, 2'd0 }; // Age: 57, HR: 98, Class: 0
mem[527] = { 8'd58, 8'd65, 2'd0 }; // Age: 58, HR: 165, Class: 0
mem[528] = { 8'd71, 8'd15, 2'd3 }; // Age: 71, HR: 115, Class: 3
mem[529] = { 8'd75, 8'd12, 2'd3 }; // Age: 75, HR: 112, Class: 3
mem[530] = { 8'd56, 8'd33, 2'd3 }; // Age: 56, HR: 133, Class: 3
mem[531] = { 8'd47, 8'd25, 2'd0 }; // Age: 47, HR: 125, Class: 0
mem[532] = { 8'd53, 8'd20, 2'd1 }; // Age: 53, HR: 120, Class: 1
mem[533] = { 8'd41, 8'd58, 2'd1 }; // Age: 41, HR: 158, Class: 1
mem[534] = { 8'd52, 8'd28, 2'd2 }; // Age: 52, HR: 128, Class: 2
mem[535] = { 8'd49, 8'd75, 2'd1 }; // Age: 49, HR: 175, Class: 1
mem[536] = { 8'd59, 8'd31, 2'd0 }; // Age: 59, HR: 131, Class: 0
mem[537] = { 8'd63, 8'd21, 2'd1 }; // Age: 63, HR: 121, Class: 1
mem[538] = { 8'd52, 8'd61, 2'd1 }; // Age: 52, HR: 161, Class: 1
mem[539] = { 8'd53, 8'd20, 2'd0 }; // Age: 53, HR: 120, Class: 0
mem[540] = { 8'd35, 8'd82, 2'd0 }; // Age: 35, HR: 182, Class: 0
mem[541] = { 8'd48, 8'd8, 2'd1 }; // Age: 48, HR: 108, Class: 1
mem[542] = { 8'd38, 8'd66, 2'd2 }; // Age: 38, HR: 166, Class: 2
mem[543] = { 8'd61, 8'd15, 2'd0 }; // Age: 61, HR: 115, Class: 0
mem[544] = { 8'd56, 8'd3, 2'd2 }; // Age: 56, HR: 103, Class: 2
mem[545] = { 8'd66, 8'd38, 2'd0 }; // Age: 66, HR: 138, Class: 0
mem[546] = { 8'd54, 8'd95, 2'd1 }; // Age: 54, HR: 195, Class: 1
mem[547] = { 8'd65, 8'd249, 2'd1 }; // Age: 65, HR: 93, Class: 1
mem[548] = { 8'd54, 8'd40, 2'd0 }; // Age: 54, HR: 140, Class: 0
mem[549] = { 8'd66, 8'd250, 2'd1 }; // Age: 66, HR: 94, Class: 1
mem[550] = { 8'd62, 8'd12, 2'd1 }; // Age: 62, HR: 112, Class: 1
mem[551] = { 8'd62, 8'd38, 2'd1 }; // Age: 62, HR: 138, Class: 1
mem[552] = { 8'd58, 8'd56, 2'd2 }; // Age: 58, HR: 156, Class: 2
mem[553] = { 8'd65, 8'd51, 2'd0 }; // Age: 65, HR: 151, Class: 0
mem[554] = { 8'd55, 8'd45, 2'd3 }; // Age: 55, HR: 145, Class: 3
mem[555] = { 8'd56, 8'd0, 2'd2 }; // Age: 56, HR: 100, Class: 2
mem[556] = { 8'd53, 8'd42, 2'd0 }; // Age: 53, HR: 142, Class: 0
mem[557] = { 8'd44, 8'd80, 2'd0 }; // Age: 44, HR: 180, Class: 0
mem[558] = { 8'd63, 8'd49, 2'd2 }; // Age: 63, HR: 149, Class: 2
mem[559] = { 8'd61, 8'd61, 2'd2 }; // Age: 61, HR: 161, Class: 2
mem[560] = { 8'd59, 8'd82, 2'd0 }; // Age: 59, HR: 182, Class: 0
mem[561] = { 8'd59, 8'd40, 2'd2 }; // Age: 59, HR: 140, Class: 2
mem[562] = { 8'd51, 8'd23, 2'd0 }; // Age: 51, HR: 123, Class: 0
mem[563] = { 8'd44, 8'd75, 2'd0 }; // Age: 44, HR: 175, Class: 0
mem[564] = { 8'd60, 8'd33, 2'd0 }; // Age: 60, HR: 133, Class: 0
mem[565] = { 8'd54, 8'd10, 2'd0 }; // Age: 54, HR: 110, Class: 0
mem[566] = { 8'd64, 8'd33, 2'd0 }; // Age: 64, HR: 133, Class: 0
mem[567] = { 8'd46, 8'd52, 2'd0 }; // Age: 46, HR: 152, Class: 0
mem[568] = { 8'd57, 8'd254, 2'd0 }; // Age: 57, HR: 98, Class: 0
mem[569] = { 8'd52, 8'd65, 2'd0 }; // Age: 52, HR: 165, Class: 0
mem[570] = { 8'd39, 8'd60, 2'd0 }; // Age: 39, HR: 160, Class: 0
mem[571] = { 8'd57, 8'd248, 2'd1 }; // Age: 57, HR: 92, Class: 1
mem[572] = { 8'd43, 8'd45, 2'd3 }; // Age: 43, HR: 145, Class: 3
mem[573] = { 8'd56, 8'd63, 2'd0 }; // Age: 56, HR: 163, Class: 0
mem[574] = { 8'd51, 8'd57, 2'd0 }; // Age: 51, HR: 157, Class: 0
mem[575] = { 8'd63, 8'd240, 2'd3 }; // Age: 63, HR: 84, Class: 3
mem[576] = { 8'd42, 8'd50, 2'd0 }; // Age: 42, HR: 150, Class: 0
mem[577] = { 8'd58, 8'd60, 2'd1 }; // Age: 58, HR: 160, Class: 1
mem[578] = { 8'd62, 8'd253, 2'd2 }; // Age: 62, HR: 97, Class: 2
mem[579] = { 8'd57, 8'd45, 2'd1 }; // Age: 57, HR: 145, Class: 1
mem[580] = { 8'd51, 8'd7, 2'd0 }; // Age: 51, HR: 107, Class: 0
mem[581] = { 8'd57, 8'd19, 2'd3 }; // Age: 57, HR: 119, Class: 3
mem[582] = { 8'd48, 8'd86, 2'd0 }; // Age: 48, HR: 186, Class: 0
mem[583] = { 8'd63, 8'd21, 2'd1 }; // Age: 63, HR: 121, Class: 1
mem[584] = { 8'd53, 8'd73, 2'd0 }; // Age: 53, HR: 173, Class: 0
mem[585] = { 8'd39, 8'd79, 2'd0 }; // Age: 39, HR: 179, Class: 0
mem[586] = { 8'd62, 8'd253, 2'd2 }; // Age: 62, HR: 97, Class: 2
mem[587] = { 8'd56, 8'd21, 2'd1 }; // Age: 56, HR: 121, Class: 1
mem[588] = { 8'd53, 8'd55, 2'd0 }; // Age: 53, HR: 155, Class: 0
mem[589] = { 8'd41, 8'd76, 2'd2 }; // Age: 41, HR: 176, Class: 2
mem[590] = { 8'd57, 8'd48, 2'd1 }; // Age: 57, HR: 148, Class: 1
mem[591] = { 8'd37, 8'd42, 2'd0 }; // Age: 37, HR: 142, Class: 0
mem[592] = { 8'd50, 8'd50, 2'd1 }; // Age: 50, HR: 150, Class: 1
mem[593] = { 8'd57, 8'd74, 2'd0 }; // Age: 57, HR: 174, Class: 0
mem[594] = { 8'd40, 8'd236, 2'd0 }; // Age: 40, HR: 80, Class: 0
mem[595] = { 8'd39, 8'd60, 2'd0 }; // Age: 39, HR: 160, Class: 0
mem[596] = { 8'd59, 8'd28, 2'd2 }; // Age: 59, HR: 128, Class: 2
mem[597] = { 8'd76, 8'd16, 2'd0 }; // Age: 76, HR: 116, Class: 0
mem[598] = { 8'd38, 8'd66, 2'd1 }; // Age: 38, HR: 166, Class: 1
mem[599] = { 8'd68, 8'd51, 2'd0 }; // Age: 68, HR: 151, Class: 0
mem[600] = { 8'd57, 8'd26, 2'd0 }; // Age: 57, HR: 126, Class: 0
mem[601] = { 8'd56, 8'd254, 2'd1 }; // Age: 56, HR: 98, Class: 1
mem[602] = { 8'd57, 8'd254, 2'd2 }; // Age: 57, HR: 98, Class: 2
mem[603] = { 8'd62, 8'd23, 2'd1 }; // Age: 62, HR: 123, Class: 1
mem[604] = { 8'd60, 8'd10, 2'd3 }; // Age: 60, HR: 110, Class: 3
mem[605] = { 8'd45, 8'd40, 2'd0 }; // Age: 45, HR: 140, Class: 0
mem[606] = { 8'd54, 8'd247, 2'd1 }; // Age: 54, HR: 91, Class: 1
mem[607] = { 8'd62, 8'd34, 2'd1 }; // Age: 62, HR: 134, Class: 1
mem[608] = { 8'd52, 8'd40, 2'd0 }; // Age: 52, HR: 140, Class: 0
mem[609] = { 8'd43, 8'd40, 2'd2 }; // Age: 43, HR: 140, Class: 2
mem[610] = { 8'd59, 8'd34, 2'd2 }; // Age: 59, HR: 134, Class: 2
mem[611] = { 8'd72, 8'd30, 2'd2 }; // Age: 72, HR: 130, Class: 2
mem[612] = { 8'd58, 8'd255, 2'd1 }; // Age: 58, HR: 99, Class: 1
mem[613] = { 8'd50, 8'd35, 2'd0 }; // Age: 50, HR: 135, Class: 0
mem[614] = { 8'd54, 8'd59, 2'd0 }; // Age: 54, HR: 159, Class: 0
mem[615] = { 8'd37, 8'd65, 2'd0 }; // Age: 37, HR: 165, Class: 0
mem[616] = { 8'd71, 8'd62, 2'd0 }; // Age: 71, HR: 162, Class: 0
mem[617] = { 8'd44, 8'd50, 2'd1 }; // Age: 44, HR: 150, Class: 1
mem[618] = { 8'd61, 8'd61, 2'd2 }; // Age: 61, HR: 161, Class: 2
mem[619] = { 8'd48, 8'd75, 2'd0 }; // Age: 48, HR: 175, Class: 0
mem[620] = { 8'd56, 8'd53, 2'd0 }; // Age: 56, HR: 153, Class: 0
mem[621] = { 8'd40, 8'd44, 2'd2 }; // Age: 40, HR: 144, Class: 2
mem[622] = { 8'd57, 8'd74, 2'd1 }; // Age: 57, HR: 174, Class: 1
mem[623] = { 8'd64, 8'd5, 2'd0 }; // Age: 64, HR: 105, Class: 0
mem[624] = { 8'd38, 8'd34, 2'd1 }; // Age: 38, HR: 134, Class: 1
mem[625] = { 8'd61, 8'd242, 2'd3 }; // Age: 61, HR: 86, Class: 3
mem[626] = { 8'd44, 8'd79, 2'd0 }; // Age: 44, HR: 179, Class: 0
mem[627] = { 8'd60, 8'd41, 2'd3 }; // Age: 60, HR: 141, Class: 3
mem[628] = { 8'd60, 8'd40, 2'd1 }; // Age: 60, HR: 140, Class: 1
mem[629] = { 8'd51, 8'd49, 2'd0 }; // Age: 51, HR: 149, Class: 0
mem[630] = { 8'd57, 8'd44, 2'd2 }; // Age: 57, HR: 144, Class: 2
mem[631] = { 8'd38, 8'd50, 2'd2 }; // Age: 38, HR: 150, Class: 2
mem[632] = { 8'd38, 8'd56, 2'd1 }; // Age: 38, HR: 156, Class: 1
mem[633] = { 8'd50, 8'd40, 2'd0 }; // Age: 50, HR: 140, Class: 0
mem[634] = { 8'd62, 8'd253, 2'd2 }; // Age: 62, HR: 97, Class: 2
mem[635] = { 8'd47, 8'd20, 2'd1 }; // Age: 47, HR: 120, Class: 1
mem[636] = { 8'd67, 8'd25, 2'd3 }; // Age: 67, HR: 125, Class: 3
mem[637] = { 8'd64, 8'd2, 2'd3 }; // Age: 64, HR: 102, Class: 3
mem[638] = { 8'd41, 8'd70, 2'd1 }; // Age: 41, HR: 170, Class: 1
mem[639] = { 8'd51, 8'd27, 2'd2 }; // Age: 51, HR: 127, Class: 2
mem[640] = { 8'd34, 8'd80, 2'd1 }; // Age: 34, HR: 180, Class: 1
mem[641] = { 8'd44, 8'd77, 2'd1 }; // Age: 44, HR: 177, Class: 1
mem[642] = { 8'd50, 8'd10, 2'd0 }; // Age: 50, HR: 110, Class: 0
mem[643] = { 8'd45, 8'd80, 2'd0 }; // Age: 45, HR: 180, Class: 0
mem[644] = { 8'd51, 8'd20, 2'd0 }; // Age: 51, HR: 120, Class: 0
mem[645] = { 8'd56, 8'd40, 2'd0 }; // Age: 56, HR: 140, Class: 0
mem[646] = { 8'd66, 8'd52, 2'd0 }; // Age: 66, HR: 152, Class: 0
mem[647] = { 8'd55, 8'd25, 2'd1 }; // Age: 55, HR: 125, Class: 1
mem[648] = { 8'd60, 8'd30, 2'd1 }; // Age: 60, HR: 130, Class: 1
mem[649] = { 8'd48, 8'd48, 2'd0 }; // Age: 48, HR: 148, Class: 0
mem[650] = { 8'd54, 8'd22, 2'd0 }; // Age: 54, HR: 122, Class: 0
mem[651] = { 8'd51, 8'd22, 2'd3 }; // Age: 51, HR: 122, Class: 3
mem[652] = { 8'd64, 8'd6, 2'd1 }; // Age: 64, HR: 106, Class: 1
mem[653] = { 8'd62, 8'd43, 2'd2 }; // Age: 62, HR: 143, Class: 2
mem[654] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[655] = { 8'd54, 8'd42, 2'd1 }; // Age: 54, HR: 142, Class: 1
mem[656] = { 8'd52, 8'd61, 2'd1 }; // Age: 52, HR: 161, Class: 1
mem[657] = { 8'd57, 8'd254, 2'd2 }; // Age: 57, HR: 98, Class: 2
mem[658] = { 8'd57, 8'd0, 2'd3 }; // Age: 57, HR: 100, Class: 3
mem[659] = { 8'd69, 8'd46, 2'd2 }; // Age: 69, HR: 146, Class: 2
mem[660] = { 8'd63, 8'd20, 2'd0 }; // Age: 63, HR: 120, Class: 0
mem[661] = { 8'd43, 8'd20, 2'd3 }; // Age: 43, HR: 120, Class: 3
mem[662] = { 8'd49, 8'd45, 2'd2 }; // Age: 49, HR: 145, Class: 2
mem[663] = { 8'd43, 8'd75, 2'd0 }; // Age: 43, HR: 175, Class: 0
mem[664] = { 8'd62, 8'd234, 2'd3 }; // Age: 62, HR: 78, Class: 3
mem[665] = { 8'd60, 8'd25, 2'd1 }; // Age: 60, HR: 125, Class: 1
mem[666] = { 8'd57, 8'd64, 2'd1 }; // Age: 57, HR: 164, Class: 1
mem[667] = { 8'd46, 8'd72, 2'd0 }; // Age: 46, HR: 172, Class: 0
mem[668] = { 8'd63, 8'd60, 2'd0 }; // Age: 63, HR: 160, Class: 0
mem[669] = { 8'd46, 8'd20, 2'd2 }; // Age: 46, HR: 120, Class: 2
mem[670] = { 8'd46, 8'd60, 2'd0 }; // Age: 46, HR: 160, Class: 0
mem[671] = { 8'd65, 8'd15, 2'd1 }; // Age: 65, HR: 115, Class: 1
mem[672] = { 8'd56, 8'd40, 2'd0 }; // Age: 56, HR: 140, Class: 0
mem[673] = { 8'd39, 8'd32, 2'd0 }; // Age: 39, HR: 132, Class: 0
mem[674] = { 8'd48, 8'd75, 2'd0 }; // Age: 48, HR: 175, Class: 0
mem[675] = { 8'd63, 8'd54, 2'd3 }; // Age: 63, HR: 154, Class: 3
mem[676] = { 8'd48, 8'd39, 2'd0 }; // Age: 48, HR: 139, Class: 0
mem[677] = { 8'd52, 8'd47, 2'd0 }; // Age: 52, HR: 147, Class: 0
mem[678] = { 8'd43, 8'd45, 2'd3 }; // Age: 43, HR: 145, Class: 3
mem[679] = { 8'd48, 8'd25, 2'd0 }; // Age: 48, HR: 125, Class: 0
mem[680] = { 8'd54, 8'd50, 2'd0 }; // Age: 54, HR: 150, Class: 0
mem[681] = { 8'd49, 8'd26, 2'd1 }; // Age: 49, HR: 126, Class: 1
mem[682] = { 8'd65, 8'd51, 2'd0 }; // Age: 65, HR: 151, Class: 0
mem[683] = { 8'd61, 8'd25, 2'd3 }; // Age: 61, HR: 125, Class: 3
mem[684] = { 8'd54, 8'd75, 2'd0 }; // Age: 54, HR: 175, Class: 0
mem[685] = { 8'd62, 8'd50, 2'd1 }; // Age: 62, HR: 150, Class: 1
mem[686] = { 8'd74, 8'd23, 2'd1 }; // Age: 74, HR: 123, Class: 1
mem[687] = { 8'd46, 8'd25, 2'd1 }; // Age: 46, HR: 125, Class: 1
mem[688] = { 8'd46, 8'd50, 2'd0 }; // Age: 46, HR: 150, Class: 0
mem[689] = { 8'd52, 8'd252, 2'd1 }; // Age: 52, HR: 96, Class: 1
mem[690] = { 8'd55, 8'd27, 2'd1 }; // Age: 55, HR: 127, Class: 1
mem[691] = { 8'd46, 8'd25, 2'd1 }; // Age: 46, HR: 125, Class: 1
mem[692] = { 8'd43, 8'd18, 2'd0 }; // Age: 43, HR: 118, Class: 0
mem[693] = { 8'd64, 8'd31, 2'd1 }; // Age: 64, HR: 131, Class: 1
mem[694] = { 8'd59, 8'd40, 2'd2 }; // Age: 59, HR: 140, Class: 2
mem[695] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[696] = { 8'd48, 8'd25, 2'd0 }; // Age: 48, HR: 125, Class: 0
mem[697] = { 8'd60, 8'd32, 2'd3 }; // Age: 60, HR: 132, Class: 3
mem[698] = { 8'd56, 8'd64, 2'd0 }; // Age: 56, HR: 164, Class: 0
mem[699] = { 8'd59, 8'd0, 2'd0 }; // Age: 59, HR: 100, Class: 0
mem[700] = { 8'd52, 8'd10, 2'd1 }; // Age: 52, HR: 110, Class: 1
mem[701] = { 8'd52, 8'd78, 2'd0 }; // Age: 52, HR: 178, Class: 0
mem[702] = { 8'd64, 8'd31, 2'd1 }; // Age: 64, HR: 131, Class: 1
mem[703] = { 8'd53, 8'd20, 2'd1 }; // Age: 53, HR: 120, Class: 1
mem[704] = { 8'd55, 8'd32, 2'd3 }; // Age: 55, HR: 132, Class: 3
mem[705] = { 8'd61, 8'd40, 2'd2 }; // Age: 61, HR: 140, Class: 2
mem[706] = { 8'd62, 8'd28, 2'd2 }; // Age: 62, HR: 128, Class: 2
mem[707] = { 8'd40, 8'd78, 2'd0 }; // Age: 40, HR: 178, Class: 0
mem[708] = { 8'd63, 8'd79, 2'd0 }; // Age: 63, HR: 179, Class: 0
mem[709] = { 8'd48, 8'd10, 2'd0 }; // Age: 48, HR: 110, Class: 0
mem[710] = { 8'd39, 8'd79, 2'd0 }; // Age: 39, HR: 179, Class: 0
mem[711] = { 8'd52, 8'd28, 2'd2 }; // Age: 52, HR: 128, Class: 2
mem[712] = { 8'd29, 8'd102, 2'd0 }; // Age: 29, HR: 202, Class: 0
mem[713] = { 8'd54, 8'd58, 2'd0 }; // Age: 54, HR: 158, Class: 0
mem[714] = { 8'd52, 8'd60, 2'd1 }; // Age: 52, HR: 160, Class: 1
mem[715] = { 8'd62, 8'd242, 2'd0 }; // Age: 62, HR: 86, Class: 0
mem[716] = { 8'd54, 8'd63, 2'd0 }; // Age: 54, HR: 163, Class: 0
mem[717] = { 8'd67, 8'd22, 2'd3 }; // Age: 67, HR: 122, Class: 3
mem[718] = { 8'd56, 8'd3, 2'd3 }; // Age: 56, HR: 103, Class: 3
mem[719] = { 8'd59, 8'd31, 2'd0 }; // Age: 59, HR: 131, Class: 0
mem[720] = { 8'd49, 8'd22, 2'd1 }; // Age: 49, HR: 122, Class: 1
mem[721] = { 8'd63, 8'd47, 2'd2 }; // Age: 63, HR: 147, Class: 2
mem[722] = { 8'd65, 8'd58, 2'd1 }; // Age: 65, HR: 158, Class: 1
mem[723] = { 8'd33, 8'd50, 2'd1 }; // Age: 33, HR: 150, Class: 1
mem[724] = { 8'd64, 8'd5, 2'd0 }; // Age: 64, HR: 105, Class: 0
mem[725] = { 8'd66, 8'd32, 2'd2 }; // Age: 66, HR: 132, Class: 2
mem[726] = { 8'd54, 8'd40, 2'd1 }; // Age: 54, HR: 140, Class: 1
mem[727] = { 8'd62, 8'd57, 2'd0 }; // Age: 62, HR: 157, Class: 0
mem[728] = { 8'd56, 8'd254, 2'd2 }; // Age: 56, HR: 98, Class: 2
mem[729] = { 8'd54, 8'd59, 2'd0 }; // Age: 54, HR: 159, Class: 0
mem[730] = { 8'd45, 8'd38, 2'd0 }; // Age: 45, HR: 138, Class: 0
mem[731] = { 8'd47, 8'd25, 2'd0 }; // Age: 47, HR: 125, Class: 0
mem[732] = { 8'd63, 8'd244, 2'd3 }; // Age: 63, HR: 88, Class: 3
mem[733] = { 8'd52, 8'd28, 2'd2 }; // Age: 52, HR: 128, Class: 2
mem[734] = { 8'd62, 8'd6, 2'd2 }; // Age: 62, HR: 106, Class: 2
mem[735] = { 8'd51, 8'd50, 2'd1 }; // Age: 51, HR: 150, Class: 1
mem[736] = { 8'd43, 8'd71, 2'd0 }; // Age: 43, HR: 171, Class: 0
mem[737] = { 8'd48, 8'd75, 2'd0 }; // Age: 48, HR: 175, Class: 0
mem[738] = { 8'd51, 8'd20, 2'd0 }; // Age: 51, HR: 120, Class: 0
mem[739] = { 8'd39, 8'd6, 2'd0 }; // Age: 39, HR: 106, Class: 0
mem[740] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[741] = { 8'd37, 8'd30, 2'd1 }; // Age: 37, HR: 130, Class: 1
mem[742] = { 8'd43, 8'd75, 2'd0 }; // Age: 43, HR: 175, Class: 0
mem[743] = { 8'd56, 8'd19, 2'd2 }; // Age: 56, HR: 119, Class: 2
mem[744] = { 8'd39, 8'd32, 2'd0 }; // Age: 39, HR: 132, Class: 0
mem[745] = { 8'd40, 8'd52, 2'd1 }; // Age: 40, HR: 152, Class: 1
mem[746] = { 8'd56, 8'd48, 2'd2 }; // Age: 56, HR: 148, Class: 2
mem[747] = { 8'd48, 8'd3, 2'd1 }; // Age: 48, HR: 103, Class: 1
mem[748] = { 8'd37, 8'd254, 2'd0 }; // Age: 37, HR: 98, Class: 0
mem[749] = { 8'd46, 8'd72, 2'd0 }; // Age: 46, HR: 172, Class: 0
mem[750] = { 8'd57, 8'd15, 2'd3 }; // Age: 57, HR: 115, Class: 3
mem[751] = { 8'd51, 8'd54, 2'd0 }; // Age: 51, HR: 154, Class: 0
mem[752] = { 8'd61, 8'd35, 2'd3 }; // Age: 61, HR: 135, Class: 3
mem[753] = { 8'd46, 8'd47, 2'd1 }; // Age: 46, HR: 147, Class: 1
mem[754] = { 8'd58, 8'd5, 2'd1 }; // Age: 58, HR: 105, Class: 1
mem[755] = { 8'd50, 8'd70, 2'd0 }; // Age: 50, HR: 170, Class: 0
mem[756] = { 8'd65, 8'd40, 2'd3 }; // Age: 65, HR: 140, Class: 3
mem[757] = { 8'd54, 8'd50, 2'd0 }; // Age: 54, HR: 150, Class: 0
mem[758] = { 8'd56, 8'd50, 2'd2 }; // Age: 56, HR: 150, Class: 2
mem[759] = { 8'd52, 8'd69, 2'd0 }; // Age: 52, HR: 169, Class: 0
mem[760] = { 8'd66, 8'd51, 2'd0 }; // Age: 66, HR: 151, Class: 0
mem[761] = { 8'd70, 8'd248, 2'd1 }; // Age: 70, HR: 92, Class: 1
mem[762] = { 8'd51, 8'd252, 2'd0 }; // Age: 51, HR: 96, Class: 0
mem[763] = { 8'd40, 8'd30, 2'd1 }; // Age: 40, HR: 130, Class: 1
mem[764] = { 8'd55, 8'd32, 2'd3 }; // Age: 55, HR: 132, Class: 3
mem[765] = { 8'd45, 8'd75, 2'd0 }; // Age: 45, HR: 175, Class: 0
mem[766] = { 8'd54, 8'd42, 2'd0 }; // Age: 54, HR: 142, Class: 0
mem[767] = { 8'd59, 8'd43, 2'd1 }; // Age: 59, HR: 143, Class: 1
mem[768] = { 8'd56, 8'd254, 2'd2 }; // Age: 56, HR: 98, Class: 2
mem[769] = { 8'd61, 8'd242, 2'd3 }; // Age: 61, HR: 86, Class: 3
mem[770] = { 8'd59, 8'd82, 2'd0 }; // Age: 59, HR: 182, Class: 0
mem[771] = { 8'd53, 8'd20, 2'd0 }; // Age: 53, HR: 120, Class: 0
mem[772] = { 8'd41, 8'd58, 2'd1 }; // Age: 41, HR: 158, Class: 1
mem[773] = { 8'd57, 8'd48, 2'd1 }; // Age: 57, HR: 148, Class: 1
mem[774] = { 8'd57, 8'd40, 2'd0 }; // Age: 57, HR: 140, Class: 0
mem[775] = { 8'd54, 8'd37, 2'd0 }; // Age: 54, HR: 137, Class: 0
mem[776] = { 8'd41, 8'd28, 2'd0 }; // Age: 41, HR: 128, Class: 0
mem[777] = { 8'd42, 8'd46, 2'd0 }; // Age: 42, HR: 146, Class: 0
mem[778] = { 8'd63, 8'd50, 2'd0 }; // Age: 63, HR: 150, Class: 0
mem[779] = { 8'd46, 8'd40, 2'd0 }; // Age: 46, HR: 140, Class: 0
mem[780] = { 8'd40, 8'd88, 2'd0 }; // Age: 40, HR: 188, Class: 0
mem[781] = { 8'd69, 8'd46, 2'd2 }; // Age: 69, HR: 146, Class: 2
mem[782] = { 8'd46, 8'd24, 2'd1 }; // Age: 46, HR: 124, Class: 1
mem[783] = { 8'd50, 8'd63, 2'd0 }; // Age: 50, HR: 163, Class: 0
mem[784] = { 8'd47, 8'd254, 2'd1 }; // Age: 47, HR: 98, Class: 1
mem[785] = { 8'd43, 8'd75, 2'd0 }; // Age: 43, HR: 175, Class: 0
mem[786] = { 8'd49, 8'd72, 2'd0 }; // Age: 49, HR: 172, Class: 0
mem[787] = { 8'd58, 8'd18, 2'd2 }; // Age: 58, HR: 118, Class: 2
mem[788] = { 8'd58, 8'd65, 2'd0 }; // Age: 58, HR: 165, Class: 0
mem[789] = { 8'd51, 8'd86, 2'd0 }; // Age: 51, HR: 186, Class: 0
mem[790] = { 8'd41, 8'd58, 2'd1 }; // Age: 41, HR: 158, Class: 1
mem[791] = { 8'd44, 8'd50, 2'd1 }; // Age: 44, HR: 150, Class: 1
mem[792] = { 8'd61, 8'd233, 2'd3 }; // Age: 61, HR: 77, Class: 3
mem[793] = { 8'd59, 8'd19, 2'd1 }; // Age: 59, HR: 119, Class: 1
mem[794] = { 8'd59, 8'd43, 2'd1 }; // Age: 59, HR: 143, Class: 1
mem[795] = { 8'd41, 8'd28, 2'd0 }; // Age: 41, HR: 128, Class: 0
mem[796] = { 8'd54, 8'd5, 2'd1 }; // Age: 54, HR: 105, Class: 1
mem[797] = { 8'd45, 8'd70, 2'd0 }; // Age: 45, HR: 170, Class: 0
mem[798] = { 8'd58, 8'd11, 2'd3 }; // Age: 58, HR: 111, Class: 3
mem[799] = { 8'd41, 8'd68, 2'd0 }; // Age: 41, HR: 168, Class: 0
mem[800] = { 8'd57, 8'd73, 2'd0 }; // Age: 57, HR: 173, Class: 0
mem[801] = { 8'd53, 8'd6, 2'd1 }; // Age: 53, HR: 106, Class: 1
mem[802] = { 8'd54, 8'd8, 2'd3 }; // Age: 54, HR: 108, Class: 3
mem[803] = { 8'd60, 8'd30, 2'd1 }; // Age: 60, HR: 130, Class: 1
mem[804] = { 8'd47, 8'd43, 2'd0 }; // Age: 47, HR: 143, Class: 0
mem[805] = { 8'd56, 8'd21, 2'd1 }; // Age: 56, HR: 121, Class: 1
mem[806] = { 8'd43, 8'd55, 2'd1 }; // Age: 43, HR: 155, Class: 1
mem[807] = { 8'd53, 8'd48, 2'd0 }; // Age: 53, HR: 148, Class: 0
mem[808] = { 8'd48, 8'd18, 2'd0 }; // Age: 48, HR: 118, Class: 0
mem[809] = { 8'd51, 8'd23, 2'd0 }; // Age: 51, HR: 123, Class: 0
mem[810] = { 8'd49, 8'd26, 2'd1 }; // Age: 49, HR: 126, Class: 1
mem[811] = { 8'd29, 8'd60, 2'd0 }; // Age: 29, HR: 160, Class: 0
mem[812] = { 8'd63, 8'd15, 2'd1 }; // Age: 63, HR: 115, Class: 1
mem[813] = { 8'd52, 8'd84, 2'd0 }; // Age: 52, HR: 184, Class: 0
mem[814] = { 8'd50, 8'd70, 2'd0 }; // Age: 50, HR: 170, Class: 0
mem[815] = { 8'd49, 8'd75, 2'd1 }; // Age: 49, HR: 175, Class: 1
mem[816] = { 8'd44, 8'd35, 2'd0 }; // Age: 44, HR: 135, Class: 0
mem[817] = { 8'd52, 8'd24, 2'd1 }; // Age: 52, HR: 124, Class: 1
mem[818] = { 8'd70, 8'd43, 2'd0 }; // Age: 70, HR: 143, Class: 0
mem[819] = { 8'd56, 8'd0, 2'd2 }; // Age: 56, HR: 100, Class: 2
mem[820] = { 8'd56, 8'd14, 2'd0 }; // Age: 56, HR: 114, Class: 0
mem[821] = { 8'd56, 8'd53, 2'd0 }; // Age: 56, HR: 153, Class: 0
mem[822] = { 8'd37, 8'd58, 2'd0 }; // Age: 37, HR: 158, Class: 0
mem[823] = { 8'd63, 8'd20, 2'd0 }; // Age: 63, HR: 120, Class: 0
mem[824] = { 8'd61, 8'd48, 2'd2 }; // Age: 61, HR: 148, Class: 2
mem[825] = { 8'd42, 8'd55, 2'd0 }; // Age: 42, HR: 155, Class: 0
mem[826] = { 8'd49, 8'd74, 2'd0 }; // Age: 49, HR: 174, Class: 0
mem[827] = { 8'd58, 8'd5, 2'd1 }; // Age: 58, HR: 105, Class: 1
mem[828] = { 8'd44, 8'd35, 2'd0 }; // Age: 44, HR: 135, Class: 0
mem[829] = { 8'd57, 8'd63, 2'd0 }; // Age: 57, HR: 163, Class: 0
mem[830] = { 8'd63, 8'd54, 2'd3 }; // Age: 63, HR: 154, Class: 3
mem[831] = { 8'd40, 8'd88, 2'd0 }; // Age: 40, HR: 188, Class: 0
mem[832] = { 8'd60, 8'd30, 2'd1 }; // Age: 60, HR: 130, Class: 1
mem[833] = { 8'd51, 8'd49, 2'd0 }; // Age: 51, HR: 149, Class: 0
mem[834] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[835] = { 8'd63, 8'd242, 2'd3 }; // Age: 63, HR: 86, Class: 3
mem[836] = { 8'd35, 8'd85, 2'd0 }; // Age: 35, HR: 185, Class: 0
mem[837] = { 8'd56, 8'd5, 2'd1 }; // Age: 56, HR: 105, Class: 1
mem[838] = { 8'd50, 8'd21, 2'd1 }; // Age: 50, HR: 121, Class: 1
mem[839] = { 8'd57, 8'd48, 2'd1 }; // Age: 57, HR: 148, Class: 1
mem[840] = { 8'd65, 8'd14, 2'd3 }; // Age: 65, HR: 114, Class: 3
mem[841] = { 8'd63, 8'd11, 2'd3 }; // Age: 63, HR: 111, Class: 3
mem[842] = { 8'd65, 8'd249, 2'd1 }; // Age: 65, HR: 93, Class: 1
mem[843] = { 8'd41, 8'd38, 2'd1 }; // Age: 41, HR: 138, Class: 1
mem[844] = { 8'd58, 8'd54, 2'd0 }; // Age: 58, HR: 154, Class: 0
mem[845] = { 8'd50, 8'd59, 2'd0 }; // Age: 50, HR: 159, Class: 0
mem[846] = { 8'd66, 8'd20, 2'd0 }; // Age: 66, HR: 120, Class: 0
mem[847] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[848] = { 8'd57, 8'd48, 2'd1 }; // Age: 57, HR: 148, Class: 1
mem[849] = { 8'd61, 8'd236, 2'd3 }; // Age: 61, HR: 80, Class: 3
mem[850] = { 8'd46, 8'd75, 2'd1 }; // Age: 46, HR: 175, Class: 1
mem[851] = { 8'd54, 8'd18, 2'd1 }; // Age: 54, HR: 118, Class: 1
mem[852] = { 8'd64, 8'd5, 2'd0 }; // Age: 64, HR: 105, Class: 0
mem[853] = { 8'd47, 8'd45, 2'd0 }; // Age: 47, HR: 145, Class: 0
mem[854] = { 8'd56, 8'd50, 2'd1 }; // Age: 56, HR: 150, Class: 1
mem[855] = { 8'd42, 8'd73, 2'd0 }; // Age: 42, HR: 173, Class: 0
mem[856] = { 8'd66, 8'd8, 2'd3 }; // Age: 66, HR: 108, Class: 3
mem[857] = { 8'd54, 8'd5, 2'd1 }; // Age: 54, HR: 105, Class: 1
mem[858] = { 8'd54, 8'd37, 2'd0 }; // Age: 54, HR: 137, Class: 0
mem[859] = { 8'd53, 8'd55, 2'd1 }; // Age: 53, HR: 155, Class: 1
mem[860] = { 8'd58, 8'd18, 2'd2 }; // Age: 58, HR: 118, Class: 2
mem[861] = { 8'd63, 8'd60, 2'd0 }; // Age: 63, HR: 160, Class: 0
mem[862] = { 8'd41, 8'd63, 2'd0 }; // Age: 41, HR: 163, Class: 0
mem[863] = { 8'd57, 8'd26, 2'd0 }; // Age: 57, HR: 126, Class: 0
mem[864] = { 8'd41, 8'd72, 2'd0 }; // Age: 41, HR: 172, Class: 0
mem[865] = { 8'd63, 8'd32, 2'd3 }; // Age: 63, HR: 132, Class: 3
mem[866] = { 8'd48, 8'd10, 2'd1 }; // Age: 48, HR: 110, Class: 1
mem[867] = { 8'd44, 8'd70, 2'd0 }; // Age: 44, HR: 170, Class: 0
mem[868] = { 8'd54, 8'd13, 2'd2 }; // Age: 54, HR: 113, Class: 2
mem[869] = { 8'd47, 8'd52, 2'd1 }; // Age: 47, HR: 152, Class: 1
mem[870] = { 8'd53, 8'd251, 2'd3 }; // Age: 53, HR: 95, Class: 3
mem[871] = { 8'd49, 8'd62, 2'd0 }; // Age: 49, HR: 162, Class: 0
mem[872] = { 8'd52, 8'd47, 2'd0 }; // Age: 52, HR: 147, Class: 0
mem[873] = { 8'd75, 8'd8, 2'd1 }; // Age: 75, HR: 108, Class: 1
mem[874] = { 8'd57, 8'd252, 2'd0 }; // Age: 57, HR: 96, Class: 0
mem[875] = { 8'd47, 8'd79, 2'd0 }; // Age: 47, HR: 179, Class: 0
mem[876] = { 8'd58, 8'd31, 2'd1 }; // Age: 58, HR: 131, Class: 1
mem[877] = { 8'd46, 8'd72, 2'd0 }; // Age: 46, HR: 172, Class: 0
mem[878] = { 8'd61, 8'd254, 2'd3 }; // Age: 61, HR: 98, Class: 3
mem[879] = { 8'd59, 8'd54, 2'd0 }; // Age: 59, HR: 154, Class: 0
mem[880] = { 8'd63, 8'd244, 2'd3 }; // Age: 63, HR: 88, Class: 3
mem[881] = { 8'd62, 8'd43, 2'd2 }; // Age: 62, HR: 143, Class: 2
mem[882] = { 8'd55, 8'd50, 2'd0 }; // Age: 55, HR: 150, Class: 0
mem[883] = { 8'd42, 8'd255, 2'd2 }; // Age: 42, HR: 99, Class: 2
mem[884] = { 8'd49, 8'd39, 2'd3 }; // Age: 49, HR: 139, Class: 3
mem[885] = { 8'd52, 8'd58, 2'd0 }; // Age: 52, HR: 158, Class: 0
mem[886] = { 8'd48, 8'd3, 2'd1 }; // Age: 48, HR: 103, Class: 1
mem[887] = { 8'd46, 8'd16, 2'd0 }; // Age: 46, HR: 116, Class: 0
mem[888] = { 8'd49, 8'd60, 2'd0 }; // Age: 49, HR: 160, Class: 0
mem[889] = { 8'd53, 8'd60, 2'd0 }; // Age: 53, HR: 160, Class: 0
mem[890] = { 8'd52, 8'd20, 2'd1 }; // Age: 52, HR: 120, Class: 1
mem[891] = { 8'd57, 8'd40, 2'd0 }; // Age: 57, HR: 140, Class: 0
mem[892] = { 8'd66, 8'd8, 2'd3 }; // Age: 66, HR: 108, Class: 3
mem[893] = { 8'd54, 8'd54, 2'd1 }; // Age: 54, HR: 154, Class: 1
mem[894] = { 8'd54, 8'd55, 2'd2 }; // Age: 54, HR: 155, Class: 2
mem[895] = { 8'd58, 8'd10, 2'd2 }; // Age: 58, HR: 110, Class: 2
mem[896] = { 8'd53, 8'd32, 2'd0 }; // Age: 53, HR: 132, Class: 0
mem[897] = { 8'd58, 8'd60, 2'd1 }; // Age: 58, HR: 160, Class: 1
mem[898] = { 8'd52, 8'd10, 2'd1 }; // Age: 52, HR: 110, Class: 1
mem[899] = { 8'd60, 8'd219, 2'd3 }; // Age: 60, HR: 63, Class: 3
mem[900] = { 8'd70, 8'd248, 2'd1 }; // Age: 70, HR: 92, Class: 1
mem[901] = { 8'd54, 8'd34, 2'd0 }; // Age: 54, HR: 134, Class: 0
mem[902] = { 8'd39, 8'd82, 2'd0 }; // Age: 39, HR: 182, Class: 0
mem[903] = { 8'd58, 8'd54, 2'd0 }; // Age: 58, HR: 154, Class: 0
mem[904] = { 8'd52, 8'd72, 2'd0 }; // Age: 52, HR: 172, Class: 0
mem[905] = { 8'd51, 8'd42, 2'd0 }; // Age: 51, HR: 142, Class: 0
mem[906] = { 8'd54, 8'd22, 2'd0 }; // Age: 54, HR: 122, Class: 0
mem[907] = { 8'd63, 8'd50, 2'd0 }; // Age: 63, HR: 150, Class: 0
mem[908] = { 8'd41, 8'd68, 2'd0 }; // Age: 41, HR: 168, Class: 0
mem[909] = { 8'd61, 8'd233, 2'd3 }; // Age: 61, HR: 77, Class: 3
mem[910] = { 8'd73, 8'd21, 2'd1 }; // Age: 73, HR: 121, Class: 1
mem[911] = { 8'd69, 8'd18, 2'd2 }; // Age: 69, HR: 118, Class: 2
mem[912] = { 8'd54, 8'd55, 2'd0 }; // Age: 54, HR: 155, Class: 0
mem[913] = { 8'd54, 8'd30, 2'd0 }; // Age: 54, HR: 130, Class: 0
mem[914] = { 8'd61, 8'd15, 2'd0 }; // Age: 61, HR: 115, Class: 0
mem[915] = { 8'd65, 8'd20, 2'd3 }; // Age: 65, HR: 120, Class: 3
mem[916] = { 8'd59, 8'd61, 2'd0 }; // Age: 59, HR: 161, Class: 0
mem[917] = { 8'd40, 8'd88, 2'd0 }; // Age: 40, HR: 188, Class: 0
mem[918] = { 8'd63, 8'd72, 2'd0 }; // Age: 63, HR: 172, Class: 0
mem[919] = { 8'd67, 8'd63, 2'd3 }; // Age: 67, HR: 163, Class: 3
mem[920] = { 8'd57, 8'd248, 2'd1 }; // Age: 57, HR: 92, Class: 1
mem[921] = { 8'd55, 8'd45, 2'd3 }; // Age: 55, HR: 145, Class: 3
mem[922] = { 8'd62, 8'd40, 2'd0 }; // Age: 62, HR: 140, Class: 0
mem[923] = { 8'd60, 8'd43, 2'd1 }; // Age: 60, HR: 143, Class: 1
mem[924] = { 8'd53, 8'd62, 2'd0 }; // Age: 53, HR: 162, Class: 0
mem[925] = { 8'd35, 8'd82, 2'd0 }; // Age: 35, HR: 182, Class: 0
mem[926] = { 8'd58, 8'd10, 2'd2 }; // Age: 58, HR: 110, Class: 2
mem[927] = { 8'd29, 8'd70, 2'd0 }; // Age: 29, HR: 170, Class: 0
mem[928] = { 8'd59, 8'd34, 2'd2 }; // Age: 59, HR: 134, Class: 2
mem[929] = { 8'd44, 8'd88, 2'd0 }; // Age: 44, HR: 188, Class: 0
mem[930] = { 8'd54, 8'd16, 2'd3 }; // Age: 54, HR: 116, Class: 3
mem[931] = { 8'd47, 8'd35, 2'd0 }; // Age: 47, HR: 135, Class: 0
mem[932] = { 8'd63, 8'd240, 2'd3 }; // Age: 63, HR: 84, Class: 3
mem[933] = { 8'd56, 8'd61, 2'd0 }; // Age: 56, HR: 161, Class: 0
mem[934] = { 8'd75, 8'd12, 2'd0 }; // Age: 75, HR: 112, Class: 0
mem[935] = { 8'd48, 8'd60, 2'd0 }; // Age: 48, HR: 160, Class: 0
mem[936] = { 8'd50, 8'd56, 2'd3 }; // Age: 50, HR: 156, Class: 3
mem[937] = { 8'd59, 8'd20, 2'd1 }; // Age: 59, HR: 120, Class: 1
mem[938] = { 8'd38, 8'd73, 2'd0 }; // Age: 38, HR: 173, Class: 0
mem[939] = { 8'd58, 8'd30, 2'd3 }; // Age: 58, HR: 130, Class: 3
mem[940] = { 8'd54, 8'd8, 2'd3 }; // Age: 54, HR: 108, Class: 3
mem[941] = { 8'd57, 8'd252, 2'd0 }; // Age: 57, HR: 96, Class: 0
mem[942] = { 8'd59, 8'd25, 2'd1 }; // Age: 59, HR: 125, Class: 1
mem[943] = { 8'd44, 8'd77, 2'd1 }; // Age: 44, HR: 177, Class: 1
mem[944] = { 8'd53, 8'd42, 2'd0 }; // Age: 53, HR: 142, Class: 0
mem[945] = { 8'd57, 8'd59, 2'd0 }; // Age: 57, HR: 159, Class: 0
mem[946] = { 8'd51, 8'd20, 2'd0 }; // Age: 51, HR: 120, Class: 0
mem[947] = { 8'd65, 8'd249, 2'd1 }; // Age: 65, HR: 93, Class: 1
mem[948] = { 8'd53, 8'd6, 2'd1 }; // Age: 53, HR: 106, Class: 1
mem[949] = { 8'd58, 8'd24, 2'd2 }; // Age: 58, HR: 124, Class: 2
mem[950] = { 8'd59, 8'd17, 2'd1 }; // Age: 59, HR: 117, Class: 1
mem[951] = { 8'd29, 8'd70, 2'd0 }; // Age: 29, HR: 170, Class: 0
mem[952] = { 8'd60, 8'd57, 2'd3 }; // Age: 60, HR: 157, Class: 3
mem[953] = { 8'd57, 8'd0, 2'd1 }; // Age: 57, HR: 100, Class: 1
mem[954] = { 8'd63, 8'd60, 2'd0 }; // Age: 63, HR: 160, Class: 0
mem[955] = { 8'd39, 8'd46, 2'd0 }; // Age: 39, HR: 146, Class: 0
mem[956] = { 8'd62, 8'd8, 2'd3 }; // Age: 62, HR: 108, Class: 3
mem[957] = { 8'd53, 8'd42, 2'd0 }; // Age: 53, HR: 142, Class: 0
mem[958] = { 8'd54, 8'd40, 2'd0 }; // Age: 54, HR: 140, Class: 0
mem[959] = { 8'd31, 8'd50, 2'd0 }; // Age: 31, HR: 150, Class: 0
mem[960] = { 8'd52, 8'd68, 2'd3 }; // Age: 52, HR: 168, Class: 3
mem[961] = { 8'd57, 8'd68, 2'd0 }; // Age: 57, HR: 168, Class: 0
mem[962] = { 8'd59, 8'd24, 2'd0 }; // Age: 59, HR: 124, Class: 0
mem[963] = { 8'd39, 8'd46, 2'd0 }; // Age: 39, HR: 146, Class: 0
mem[964] = { 8'd52, 8'd26, 2'd1 }; // Age: 52, HR: 126, Class: 1
mem[965] = { 8'd59, 8'd28, 2'd2 }; // Age: 59, HR: 128, Class: 2
mem[966] = { 8'd54, 8'd56, 2'd0 }; // Age: 54, HR: 156, Class: 0
mem[967] = { 8'd51, 8'd50, 2'd1 }; // Age: 51, HR: 150, Class: 1
mem[968] = { 8'd45, 8'd48, 2'd0 }; // Age: 45, HR: 148, Class: 0
mem[969] = { 8'd29, 8'd102, 2'd0 }; // Age: 29, HR: 202, Class: 0
mem[970] = { 8'd43, 8'd20, 2'd1 }; // Age: 43, HR: 120, Class: 1
mem[971] = { 8'd62, 8'd3, 2'd3 }; // Age: 62, HR: 103, Class: 3
mem[972] = { 8'd59, 8'd45, 2'd0 }; // Age: 59, HR: 145, Class: 0
mem[973] = { 8'd48, 8'd60, 2'd0 }; // Age: 48, HR: 160, Class: 0
mem[974] = { 8'd37, 8'd58, 2'd0 }; // Age: 37, HR: 158, Class: 0
mem[975] = { 8'd67, 8'd30, 2'd2 }; // Age: 67, HR: 130, Class: 2
mem[976] = { 8'd47, 8'd254, 2'd1 }; // Age: 47, HR: 98, Class: 1
mem[977] = { 8'd56, 8'd254, 2'd1 }; // Age: 56, HR: 98, Class: 1
mem[978] = { 8'd59, 8'd40, 2'd2 }; // Age: 59, HR: 140, Class: 2
mem[979] = { 8'd54, 8'd25, 2'd1 }; // Age: 54, HR: 125, Class: 1
mem[980] = { 8'd58, 8'd6, 2'd1 }; // Age: 58, HR: 106, Class: 1
mem[981] = { 8'd44, 8'd53, 2'd2 }; // Age: 44, HR: 153, Class: 2
mem[982] = { 8'd54, 8'd37, 2'd0 }; // Age: 54, HR: 137, Class: 0
mem[983] = { 8'd43, 8'd61, 2'd0 }; // Age: 43, HR: 161, Class: 0
mem[984] = { 8'd45, 8'd75, 2'd0 }; // Age: 45, HR: 175, Class: 0
mem[985] = { 8'd55, 8'd55, 2'd3 }; // Age: 55, HR: 155, Class: 3
mem[986] = { 8'd71, 8'd62, 2'd0 }; // Age: 71, HR: 162, Class: 0
mem[987] = { 8'd61, 8'd236, 2'd3 }; // Age: 61, HR: 80, Class: 3
mem[988] = { 8'd61, 8'd46, 2'd1 }; // Age: 61, HR: 146, Class: 1
mem[989] = { 8'd55, 8'd25, 2'd1 }; // Age: 55, HR: 125, Class: 1
mem[990] = { 8'd57, 8'd0, 2'd3 }; // Age: 57, HR: 100, Class: 3
mem[991] = { 8'd42, 8'd78, 2'd0 }; // Age: 42, HR: 178, Class: 0
mem[992] = { 8'd58, 8'd13, 2'd3 }; // Age: 58, HR: 113, Class: 3
mem[993] = { 8'd63, 8'd72, 2'd0 }; // Age: 63, HR: 172, Class: 0
mem[994] = { 8'd44, 8'd70, 2'd0 }; // Age: 44, HR: 170, Class: 0
mem[995] = { 8'd54, 8'd22, 2'd1 }; // Age: 54, HR: 122, Class: 1
mem[996] = { 8'd42, 8'd52, 2'd0 }; // Age: 42, HR: 152, Class: 0
mem[997] = { 8'd63, 8'd9, 2'd1 }; // Age: 63, HR: 109, Class: 1
mem[998] = { 8'd57, 8'd43, 2'd2 }; // Age: 57, HR: 143, Class: 2
mem[999] = { 8'd68, 8'd15, 2'd0 }; // Age: 68, HR: 115, Class: 0
mem[1000] = { 8'd55, 8'd0, 2'd2 }; // Age: 55, HR: 100, Class: 2
mem[1001] = { 8'd68, 8'd15, 2'd0 }; // Age: 68, HR: 115, Class: 0
mem[1002] = { 8'd58, 8'd0, 2'd3 }; // Age: 58, HR: 100, Class: 3
mem[1003] = { 8'd62, 8'd46, 2'd0 }; // Age: 62, HR: 146, Class: 0
mem[1004] = { 8'd59, 8'd19, 2'd1 }; // Age: 59, HR: 119, Class: 1
mem[1005] = { 8'd51, 8'd42, 2'd2 }; // Age: 51, HR: 142, Class: 2
mem[1006] = { 8'd52, 8'd28, 2'd2 }; // Age: 52, HR: 128, Class: 2
mem[1007] = { 8'd41, 8'd68, 2'd0 }; // Age: 41, HR: 168, Class: 0
mem[1008] = { 8'd48, 8'd38, 2'd0 }; // Age: 48, HR: 138, Class: 0
mem[1009] = { 8'd69, 8'd40, 2'd3 }; // Age: 69, HR: 140, Class: 3
mem[1010] = { 8'd41, 8'd72, 2'd0 }; // Age: 41, HR: 172, Class: 0
mem[1011] = { 8'd55, 8'd34, 2'd0 }; // Age: 55, HR: 134, Class: 0
mem[1012] = { 8'd38, 8'd28, 2'd1 }; // Age: 38, HR: 128, Class: 1
mem[1013] = { 8'd61, 8'd13, 2'd1 }; // Age: 61, HR: 113, Class: 1
mem[1014] = { 8'd41, 8'd28, 2'd0 }; // Age: 41, HR: 128, Class: 0
mem[1015] = { 8'd46, 8'd15, 2'd1 }; // Age: 46, HR: 115, Class: 1
mem[1016] = { 8'd49, 8'd60, 2'd0 }; // Age: 49, HR: 160, Class: 0
mem[1017] = { 8'd48, 8'd59, 2'd3 }; // Age: 48, HR: 159, Class: 3
mem[1018] = { 8'd49, 8'd75, 2'd1 }; // Age: 49, HR: 175, Class: 1
mem[1019] = { 8'd54, 8'd55, 2'd2 }; // Age: 54, HR: 155, Class: 2
mem[1020] = { 8'd49, 8'd26, 2'd1 }; // Age: 49, HR: 126, Class: 1
mem[1021] = { 8'd59, 8'd30, 2'd1 }; // Age: 59, HR: 130, Class: 1
mem[1022] = { 8'd40, 8'd38, 2'd0 }; // Age: 40, HR: 138, Class: 0
mem[1023] = { 8'd58, 8'd65, 2'd3 }; // Age: 58, HR: 165, Class: 3
end

    always @(posedge clk) begin
        data_out_a <= mem[addr_a];
        data_out_b <= mem[addr_b];
    end
endmodule
